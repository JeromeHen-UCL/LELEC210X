// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"

// DATE "11/13/2024 17:08:05"

// 
// Device: Altera 10M16SAU169C8G Package UFBGA169
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module lms_dsp (
	clk_clk,
	fifo_in_wdata,
	fifo_in_wrreq,
	fifo_out_wrdata,
	fifo_out_wrreq,
	ppd_cfg_passthrough_len,
	ppd_cfg_threshold,
	ppd_cfg_clear_rs,
	ppd_cfg_enable,
	ppd_debug_count,
	ppd_debug_long_sum,
	ppd_debug_short_sum,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
input 	clk_clk;
input 	[47:0] fifo_in_wdata;
input 	fifo_in_wrreq;
output 	[47:0] fifo_out_wrdata;
output 	fifo_out_wrreq;
input 	[15:0] ppd_cfg_passthrough_len;
input 	[7:0] ppd_cfg_threshold;
input 	ppd_cfg_clear_rs;
input 	ppd_cfg_enable;
output 	[31:0] ppd_debug_count;
output 	[31:0] ppd_debug_long_sum;
output 	[31:0] ppd_debug_short_sum;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \packet_presence_detection_0|counter_inst|count_reg[0]~q ;
wire \packet_presence_detection_0|running_sum_inst|short_sum_reg[0]~q ;
wire \packet_presence_detection_0|running_sum_inst|short_sum_reg[1]~q ;
wire \packet_presence_detection_0|running_sum_inst|short_sum_reg[2]~q ;
wire \packet_presence_detection_0|running_sum_inst|short_sum_reg[3]~q ;
wire \packet_presence_detection_0|running_sum_inst|short_sum_reg[4]~q ;
wire \packet_presence_detection_0|running_sum_inst|short_sum_reg[5]~q ;
wire \packet_presence_detection_0|running_sum_inst|short_sum_reg[6]~q ;
wire \packet_presence_detection_0|running_sum_inst|short_sum_reg[7]~q ;
wire \packet_presence_detection_0|running_sum_inst|short_sum_reg[8]~q ;
wire \packet_presence_detection_0|running_sum_inst|short_sum_reg[9]~q ;
wire \packet_presence_detection_0|running_sum_inst|short_sum_reg[10]~q ;
wire \packet_presence_detection_0|running_sum_inst|short_sum_reg[11]~q ;
wire \packet_presence_detection_0|running_sum_inst|short_sum_reg[12]~q ;
wire \packet_presence_detection_0|running_sum_inst|short_sum_reg[13]~q ;
wire \packet_presence_detection_0|running_sum_inst|short_sum_reg[14]~q ;
wire \packet_presence_detection_0|running_sum_inst|short_sum_reg[15]~q ;
wire \packet_presence_detection_0|running_sum_inst|short_sum_reg[16]~q ;
wire \packet_presence_detection_0|running_sum_inst|short_sum_reg[17]~q ;
wire \avs2fifo_0|wrdata_reg[0]~q ;
wire \avs2fifo_0|wrdata_reg[1]~q ;
wire \avs2fifo_0|wrdata_reg[2]~q ;
wire \avs2fifo_0|wrdata_reg[3]~q ;
wire \avs2fifo_0|wrdata_reg[4]~q ;
wire \avs2fifo_0|wrdata_reg[5]~q ;
wire \avs2fifo_0|wrdata_reg[6]~q ;
wire \avs2fifo_0|wrdata_reg[7]~q ;
wire \avs2fifo_0|wrdata_reg[8]~q ;
wire \avs2fifo_0|wrdata_reg[9]~q ;
wire \avs2fifo_0|wrdata_reg[10]~q ;
wire \avs2fifo_0|wrdata_reg[11]~q ;
wire \avs2fifo_0|wrdata_reg[12]~q ;
wire \avs2fifo_0|wrdata_reg[13]~q ;
wire \avs2fifo_0|wrdata_reg[14]~q ;
wire \avs2fifo_0|wrdata_reg[15]~q ;
wire \avs2fifo_0|wrdata_reg[16]~q ;
wire \avs2fifo_0|wrdata_reg[17]~q ;
wire \avs2fifo_0|wrdata_reg[18]~q ;
wire \avs2fifo_0|wrdata_reg[19]~q ;
wire \avs2fifo_0|wrdata_reg[20]~q ;
wire \avs2fifo_0|wrdata_reg[21]~q ;
wire \avs2fifo_0|wrdata_reg[22]~q ;
wire \avs2fifo_0|wrdata_reg[23]~q ;
wire \avs2fifo_0|wrdata_reg[24]~q ;
wire \avs2fifo_0|wrdata_reg[25]~q ;
wire \avs2fifo_0|wrdata_reg[26]~q ;
wire \avs2fifo_0|wrdata_reg[27]~q ;
wire \avs2fifo_0|wrdata_reg[28]~q ;
wire \avs2fifo_0|wrdata_reg[29]~q ;
wire \avs2fifo_0|wrdata_reg[30]~q ;
wire \avs2fifo_0|wrdata_reg[31]~q ;
wire \avs2fifo_0|wrdata_reg[32]~q ;
wire \avs2fifo_0|wrdata_reg[33]~q ;
wire \avs2fifo_0|wrdata_reg[34]~q ;
wire \avs2fifo_0|wrdata_reg[35]~q ;
wire \avs2fifo_0|wrdata_reg[36]~q ;
wire \avs2fifo_0|wrdata_reg[37]~q ;
wire \avs2fifo_0|wrdata_reg[38]~q ;
wire \avs2fifo_0|wrdata_reg[39]~q ;
wire \avs2fifo_0|wrdata_reg[40]~q ;
wire \avs2fifo_0|wrdata_reg[41]~q ;
wire \avs2fifo_0|wrdata_reg[42]~q ;
wire \avs2fifo_0|wrdata_reg[43]~q ;
wire \avs2fifo_0|wrdata_reg[44]~q ;
wire \avs2fifo_0|wrdata_reg[45]~q ;
wire \avs2fifo_0|wrdata_reg[46]~q ;
wire \avs2fifo_0|wrdata_reg[47]~q ;
wire \avs2fifo_0|wrreq_reg~q ;
wire \packet_presence_detection_0|counter_inst|count_reg[1]~q ;
wire \packet_presence_detection_0|counter_inst|count_reg[2]~q ;
wire \packet_presence_detection_0|counter_inst|count_reg[3]~q ;
wire \packet_presence_detection_0|counter_inst|count_reg[4]~q ;
wire \packet_presence_detection_0|counter_inst|count_reg[5]~q ;
wire \packet_presence_detection_0|counter_inst|count_reg[6]~q ;
wire \packet_presence_detection_0|counter_inst|count_reg[7]~q ;
wire \packet_presence_detection_0|counter_inst|count_reg[8]~q ;
wire \packet_presence_detection_0|counter_inst|count_reg[9]~q ;
wire \packet_presence_detection_0|counter_inst|count_reg[10]~q ;
wire \packet_presence_detection_0|counter_inst|count_reg[11]~q ;
wire \packet_presence_detection_0|counter_inst|count_reg[12]~q ;
wire \packet_presence_detection_0|counter_inst|count_reg[13]~q ;
wire \packet_presence_detection_0|counter_inst|count_reg[14]~q ;
wire \packet_presence_detection_0|counter_inst|count_reg[15]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[0]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[1]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[2]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[3]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[4]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[5]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[6]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[7]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[8]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[9]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[10]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[11]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[12]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[13]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[14]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[15]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[16]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[17]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[18]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[19]~q ;
wire \packet_presence_detection_0|running_sum_inst|long_shift_rescale[20]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[0]~q ;
wire \rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[1]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[2]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[3]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[4]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[5]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[6]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[7]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[8]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[9]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[10]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[11]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[12]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[13]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[14]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[15]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[16]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[17]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[18]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[19]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[20]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[21]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[22]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[23]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[24]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[25]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[26]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[27]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[28]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[29]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[30]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[31]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[32]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[33]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[34]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[35]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[36]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[37]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[38]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[39]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[40]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[41]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[42]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[43]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[44]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[45]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[46]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_data[47]~q ;
wire \avalon_st_adapter|data_format_adapter_0|out_valid~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[12]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[0]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[11]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[10]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[9]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[8]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[7]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[6]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[5]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[4]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[3]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[2]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[1]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[23]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[22]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[21]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[20]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[19]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[18]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[17]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[16]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[15]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[14]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[13]~q ;
wire \fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_valid~q ;
wire \packet_presence_detection_0|avalon_streaming_source_data[0]~1_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[1]~2_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[2]~3_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[3]~4_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[4]~5_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[5]~6_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[6]~7_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[7]~8_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[8]~9_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[9]~10_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[10]~11_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[11]~12_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[12]~13_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[13]~14_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[14]~15_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[15]~16_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[16]~17_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[17]~18_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[18]~19_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[19]~20_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[20]~21_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[21]~22_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[22]~23_combout ;
wire \packet_presence_detection_0|avalon_streaming_source_data[23]~24_combout ;
wire \packet_presence_detection_0|delay_line_inst|delay_reg[3][24]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_valid~q ;
wire \fifo2avs_0|valid_reg~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[21]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[20]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[19]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[18]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[17]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[16]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[15]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[14]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[12]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[13]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[9]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[8]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[7]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[6]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[5]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[4]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[3]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[2]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[0]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[1]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[11]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[10]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[23]~q ;
wire \avalon_st_adapter_001|data_format_adapter_0|out_data[22]~q ;
wire \fifo2avs_0|data_reg[21]~q ;
wire \fifo2avs_0|data_reg[45]~q ;
wire \fifo2avs_0|data_reg[20]~q ;
wire \fifo2avs_0|data_reg[44]~q ;
wire \fifo2avs_0|data_reg[19]~q ;
wire \fifo2avs_0|data_reg[43]~q ;
wire \fifo2avs_0|data_reg[18]~q ;
wire \fifo2avs_0|data_reg[42]~q ;
wire \fifo2avs_0|data_reg[17]~q ;
wire \fifo2avs_0|data_reg[41]~q ;
wire \fifo2avs_0|data_reg[16]~q ;
wire \fifo2avs_0|data_reg[40]~q ;
wire \fifo2avs_0|data_reg[15]~q ;
wire \fifo2avs_0|data_reg[39]~q ;
wire \fifo2avs_0|data_reg[14]~q ;
wire \fifo2avs_0|data_reg[38]~q ;
wire \fifo2avs_0|data_reg[12]~q ;
wire \fifo2avs_0|data_reg[36]~q ;
wire \fifo2avs_0|data_reg[13]~q ;
wire \fifo2avs_0|data_reg[37]~q ;
wire \fifo2avs_0|data_reg[9]~q ;
wire \fifo2avs_0|data_reg[33]~q ;
wire \fifo2avs_0|data_reg[8]~q ;
wire \fifo2avs_0|data_reg[32]~q ;
wire \fifo2avs_0|data_reg[7]~q ;
wire \fifo2avs_0|data_reg[31]~q ;
wire \fifo2avs_0|data_reg[6]~q ;
wire \fifo2avs_0|data_reg[30]~q ;
wire \fifo2avs_0|data_reg[5]~q ;
wire \fifo2avs_0|data_reg[29]~q ;
wire \fifo2avs_0|data_reg[4]~q ;
wire \fifo2avs_0|data_reg[28]~q ;
wire \fifo2avs_0|data_reg[3]~q ;
wire \fifo2avs_0|data_reg[27]~q ;
wire \fifo2avs_0|data_reg[2]~q ;
wire \fifo2avs_0|data_reg[26]~q ;
wire \fifo2avs_0|data_reg[0]~q ;
wire \fifo2avs_0|data_reg[24]~q ;
wire \fifo2avs_0|data_reg[1]~q ;
wire \fifo2avs_0|data_reg[25]~q ;
wire \fifo2avs_0|data_reg[11]~q ;
wire \fifo2avs_0|data_reg[35]~q ;
wire \fifo2avs_0|data_reg[10]~q ;
wire \fifo2avs_0|data_reg[34]~q ;
wire \fifo2avs_0|data_reg[23]~q ;
wire \fifo2avs_0|data_reg[47]~q ;
wire \fifo2avs_0|data_reg[22]~q ;
wire \fifo2avs_0|data_reg[46]~q ;
wire \~GND~combout ;
wire \clk_clk~input_o ;
wire \ppd_cfg_passthrough_len[15]~input_o ;
wire \ppd_cfg_passthrough_len[14]~input_o ;
wire \ppd_cfg_passthrough_len[13]~input_o ;
wire \ppd_cfg_passthrough_len[12]~input_o ;
wire \ppd_cfg_passthrough_len[11]~input_o ;
wire \ppd_cfg_passthrough_len[10]~input_o ;
wire \ppd_cfg_passthrough_len[9]~input_o ;
wire \ppd_cfg_passthrough_len[8]~input_o ;
wire \ppd_cfg_passthrough_len[7]~input_o ;
wire \ppd_cfg_passthrough_len[6]~input_o ;
wire \ppd_cfg_passthrough_len[5]~input_o ;
wire \ppd_cfg_passthrough_len[4]~input_o ;
wire \ppd_cfg_passthrough_len[3]~input_o ;
wire \ppd_cfg_passthrough_len[2]~input_o ;
wire \ppd_cfg_passthrough_len[1]~input_o ;
wire \ppd_cfg_passthrough_len[0]~input_o ;
wire \ppd_cfg_clear_rs~input_o ;
wire \reset_reset_n~input_o ;
wire \ppd_cfg_threshold[0]~input_o ;
wire \ppd_cfg_threshold[1]~input_o ;
wire \ppd_cfg_threshold[2]~input_o ;
wire \ppd_cfg_threshold[3]~input_o ;
wire \ppd_cfg_threshold[4]~input_o ;
wire \ppd_cfg_threshold[5]~input_o ;
wire \ppd_cfg_threshold[6]~input_o ;
wire \ppd_cfg_threshold[7]~input_o ;
wire \ppd_cfg_enable~input_o ;
wire \fifo_in_wrreq~input_o ;
wire \fifo_in_wdata[21]~input_o ;
wire \fifo_in_wdata[45]~input_o ;
wire \fifo_in_wdata[20]~input_o ;
wire \fifo_in_wdata[44]~input_o ;
wire \fifo_in_wdata[19]~input_o ;
wire \fifo_in_wdata[43]~input_o ;
wire \fifo_in_wdata[18]~input_o ;
wire \fifo_in_wdata[42]~input_o ;
wire \fifo_in_wdata[17]~input_o ;
wire \fifo_in_wdata[41]~input_o ;
wire \fifo_in_wdata[16]~input_o ;
wire \fifo_in_wdata[40]~input_o ;
wire \fifo_in_wdata[15]~input_o ;
wire \fifo_in_wdata[39]~input_o ;
wire \fifo_in_wdata[14]~input_o ;
wire \fifo_in_wdata[38]~input_o ;
wire \fifo_in_wdata[12]~input_o ;
wire \fifo_in_wdata[36]~input_o ;
wire \fifo_in_wdata[13]~input_o ;
wire \fifo_in_wdata[37]~input_o ;
wire \fifo_in_wdata[9]~input_o ;
wire \fifo_in_wdata[33]~input_o ;
wire \fifo_in_wdata[8]~input_o ;
wire \fifo_in_wdata[32]~input_o ;
wire \fifo_in_wdata[7]~input_o ;
wire \fifo_in_wdata[31]~input_o ;
wire \fifo_in_wdata[6]~input_o ;
wire \fifo_in_wdata[30]~input_o ;
wire \fifo_in_wdata[5]~input_o ;
wire \fifo_in_wdata[29]~input_o ;
wire \fifo_in_wdata[4]~input_o ;
wire \fifo_in_wdata[28]~input_o ;
wire \fifo_in_wdata[3]~input_o ;
wire \fifo_in_wdata[27]~input_o ;
wire \fifo_in_wdata[2]~input_o ;
wire \fifo_in_wdata[26]~input_o ;
wire \fifo_in_wdata[0]~input_o ;
wire \fifo_in_wdata[24]~input_o ;
wire \fifo_in_wdata[1]~input_o ;
wire \fifo_in_wdata[25]~input_o ;
wire \fifo_in_wdata[11]~input_o ;
wire \fifo_in_wdata[35]~input_o ;
wire \fifo_in_wdata[10]~input_o ;
wire \fifo_in_wdata[34]~input_o ;
wire \fifo_in_wdata[23]~input_o ;
wire \fifo_in_wdata[47]~input_o ;
wire \fifo_in_wdata[22]~input_o ;
wire \fifo_in_wdata[46]~input_o ;


lms_dsp_altera_reset_controller rst_controller(
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk_clk(\clk_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

lms_dsp_lms_dsp_avalon_st_adapter_001 avalon_st_adapter_001(
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.out_valid(\avalon_st_adapter_001|data_format_adapter_0|out_valid~q ),
	.valid_reg(\fifo2avs_0|valid_reg~q ),
	.out_data_21(\avalon_st_adapter_001|data_format_adapter_0|out_data[21]~q ),
	.out_data_20(\avalon_st_adapter_001|data_format_adapter_0|out_data[20]~q ),
	.out_data_19(\avalon_st_adapter_001|data_format_adapter_0|out_data[19]~q ),
	.out_data_18(\avalon_st_adapter_001|data_format_adapter_0|out_data[18]~q ),
	.out_data_17(\avalon_st_adapter_001|data_format_adapter_0|out_data[17]~q ),
	.out_data_16(\avalon_st_adapter_001|data_format_adapter_0|out_data[16]~q ),
	.out_data_15(\avalon_st_adapter_001|data_format_adapter_0|out_data[15]~q ),
	.out_data_14(\avalon_st_adapter_001|data_format_adapter_0|out_data[14]~q ),
	.out_data_12(\avalon_st_adapter_001|data_format_adapter_0|out_data[12]~q ),
	.out_data_13(\avalon_st_adapter_001|data_format_adapter_0|out_data[13]~q ),
	.out_data_9(\avalon_st_adapter_001|data_format_adapter_0|out_data[9]~q ),
	.out_data_8(\avalon_st_adapter_001|data_format_adapter_0|out_data[8]~q ),
	.out_data_7(\avalon_st_adapter_001|data_format_adapter_0|out_data[7]~q ),
	.out_data_6(\avalon_st_adapter_001|data_format_adapter_0|out_data[6]~q ),
	.out_data_5(\avalon_st_adapter_001|data_format_adapter_0|out_data[5]~q ),
	.out_data_4(\avalon_st_adapter_001|data_format_adapter_0|out_data[4]~q ),
	.out_data_3(\avalon_st_adapter_001|data_format_adapter_0|out_data[3]~q ),
	.out_data_2(\avalon_st_adapter_001|data_format_adapter_0|out_data[2]~q ),
	.out_data_0(\avalon_st_adapter_001|data_format_adapter_0|out_data[0]~q ),
	.out_data_1(\avalon_st_adapter_001|data_format_adapter_0|out_data[1]~q ),
	.out_data_11(\avalon_st_adapter_001|data_format_adapter_0|out_data[11]~q ),
	.out_data_10(\avalon_st_adapter_001|data_format_adapter_0|out_data[10]~q ),
	.out_data_23(\avalon_st_adapter_001|data_format_adapter_0|out_data[23]~q ),
	.out_data_22(\avalon_st_adapter_001|data_format_adapter_0|out_data[22]~q ),
	.data_reg_21(\fifo2avs_0|data_reg[21]~q ),
	.data_reg_45(\fifo2avs_0|data_reg[45]~q ),
	.data_reg_20(\fifo2avs_0|data_reg[20]~q ),
	.data_reg_44(\fifo2avs_0|data_reg[44]~q ),
	.data_reg_19(\fifo2avs_0|data_reg[19]~q ),
	.data_reg_43(\fifo2avs_0|data_reg[43]~q ),
	.data_reg_18(\fifo2avs_0|data_reg[18]~q ),
	.data_reg_42(\fifo2avs_0|data_reg[42]~q ),
	.data_reg_17(\fifo2avs_0|data_reg[17]~q ),
	.data_reg_41(\fifo2avs_0|data_reg[41]~q ),
	.data_reg_16(\fifo2avs_0|data_reg[16]~q ),
	.data_reg_40(\fifo2avs_0|data_reg[40]~q ),
	.data_reg_15(\fifo2avs_0|data_reg[15]~q ),
	.data_reg_39(\fifo2avs_0|data_reg[39]~q ),
	.data_reg_14(\fifo2avs_0|data_reg[14]~q ),
	.data_reg_38(\fifo2avs_0|data_reg[38]~q ),
	.data_reg_12(\fifo2avs_0|data_reg[12]~q ),
	.data_reg_36(\fifo2avs_0|data_reg[36]~q ),
	.data_reg_13(\fifo2avs_0|data_reg[13]~q ),
	.data_reg_37(\fifo2avs_0|data_reg[37]~q ),
	.data_reg_9(\fifo2avs_0|data_reg[9]~q ),
	.data_reg_33(\fifo2avs_0|data_reg[33]~q ),
	.data_reg_8(\fifo2avs_0|data_reg[8]~q ),
	.data_reg_32(\fifo2avs_0|data_reg[32]~q ),
	.data_reg_7(\fifo2avs_0|data_reg[7]~q ),
	.data_reg_31(\fifo2avs_0|data_reg[31]~q ),
	.data_reg_6(\fifo2avs_0|data_reg[6]~q ),
	.data_reg_30(\fifo2avs_0|data_reg[30]~q ),
	.data_reg_5(\fifo2avs_0|data_reg[5]~q ),
	.data_reg_29(\fifo2avs_0|data_reg[29]~q ),
	.data_reg_4(\fifo2avs_0|data_reg[4]~q ),
	.data_reg_28(\fifo2avs_0|data_reg[28]~q ),
	.data_reg_3(\fifo2avs_0|data_reg[3]~q ),
	.data_reg_27(\fifo2avs_0|data_reg[27]~q ),
	.data_reg_2(\fifo2avs_0|data_reg[2]~q ),
	.data_reg_26(\fifo2avs_0|data_reg[26]~q ),
	.data_reg_0(\fifo2avs_0|data_reg[0]~q ),
	.data_reg_24(\fifo2avs_0|data_reg[24]~q ),
	.data_reg_1(\fifo2avs_0|data_reg[1]~q ),
	.data_reg_25(\fifo2avs_0|data_reg[25]~q ),
	.data_reg_11(\fifo2avs_0|data_reg[11]~q ),
	.data_reg_35(\fifo2avs_0|data_reg[35]~q ),
	.data_reg_10(\fifo2avs_0|data_reg[10]~q ),
	.data_reg_34(\fifo2avs_0|data_reg[34]~q ),
	.data_reg_23(\fifo2avs_0|data_reg[23]~q ),
	.data_reg_47(\fifo2avs_0|data_reg[47]~q ),
	.data_reg_22(\fifo2avs_0|data_reg[22]~q ),
	.data_reg_46(\fifo2avs_0|data_reg[46]~q ),
	.clk_clk(\clk_clk~input_o ));

lms_dsp_lms_dsp_avalon_st_adapter avalon_st_adapter(
	.out_data_0(\avalon_st_adapter|data_format_adapter_0|out_data[0]~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.out_data_1(\avalon_st_adapter|data_format_adapter_0|out_data[1]~q ),
	.out_data_2(\avalon_st_adapter|data_format_adapter_0|out_data[2]~q ),
	.out_data_3(\avalon_st_adapter|data_format_adapter_0|out_data[3]~q ),
	.out_data_4(\avalon_st_adapter|data_format_adapter_0|out_data[4]~q ),
	.out_data_5(\avalon_st_adapter|data_format_adapter_0|out_data[5]~q ),
	.out_data_6(\avalon_st_adapter|data_format_adapter_0|out_data[6]~q ),
	.out_data_7(\avalon_st_adapter|data_format_adapter_0|out_data[7]~q ),
	.out_data_8(\avalon_st_adapter|data_format_adapter_0|out_data[8]~q ),
	.out_data_9(\avalon_st_adapter|data_format_adapter_0|out_data[9]~q ),
	.out_data_10(\avalon_st_adapter|data_format_adapter_0|out_data[10]~q ),
	.out_data_11(\avalon_st_adapter|data_format_adapter_0|out_data[11]~q ),
	.out_data_12(\avalon_st_adapter|data_format_adapter_0|out_data[12]~q ),
	.out_data_13(\avalon_st_adapter|data_format_adapter_0|out_data[13]~q ),
	.out_data_14(\avalon_st_adapter|data_format_adapter_0|out_data[14]~q ),
	.out_data_15(\avalon_st_adapter|data_format_adapter_0|out_data[15]~q ),
	.out_data_16(\avalon_st_adapter|data_format_adapter_0|out_data[16]~q ),
	.out_data_17(\avalon_st_adapter|data_format_adapter_0|out_data[17]~q ),
	.out_data_18(\avalon_st_adapter|data_format_adapter_0|out_data[18]~q ),
	.out_data_19(\avalon_st_adapter|data_format_adapter_0|out_data[19]~q ),
	.out_data_20(\avalon_st_adapter|data_format_adapter_0|out_data[20]~q ),
	.out_data_21(\avalon_st_adapter|data_format_adapter_0|out_data[21]~q ),
	.out_data_22(\avalon_st_adapter|data_format_adapter_0|out_data[22]~q ),
	.out_data_23(\avalon_st_adapter|data_format_adapter_0|out_data[23]~q ),
	.out_data_24(\avalon_st_adapter|data_format_adapter_0|out_data[24]~q ),
	.out_data_25(\avalon_st_adapter|data_format_adapter_0|out_data[25]~q ),
	.out_data_26(\avalon_st_adapter|data_format_adapter_0|out_data[26]~q ),
	.out_data_27(\avalon_st_adapter|data_format_adapter_0|out_data[27]~q ),
	.out_data_28(\avalon_st_adapter|data_format_adapter_0|out_data[28]~q ),
	.out_data_29(\avalon_st_adapter|data_format_adapter_0|out_data[29]~q ),
	.out_data_30(\avalon_st_adapter|data_format_adapter_0|out_data[30]~q ),
	.out_data_31(\avalon_st_adapter|data_format_adapter_0|out_data[31]~q ),
	.out_data_32(\avalon_st_adapter|data_format_adapter_0|out_data[32]~q ),
	.out_data_33(\avalon_st_adapter|data_format_adapter_0|out_data[33]~q ),
	.out_data_34(\avalon_st_adapter|data_format_adapter_0|out_data[34]~q ),
	.out_data_35(\avalon_st_adapter|data_format_adapter_0|out_data[35]~q ),
	.out_data_36(\avalon_st_adapter|data_format_adapter_0|out_data[36]~q ),
	.out_data_37(\avalon_st_adapter|data_format_adapter_0|out_data[37]~q ),
	.out_data_38(\avalon_st_adapter|data_format_adapter_0|out_data[38]~q ),
	.out_data_39(\avalon_st_adapter|data_format_adapter_0|out_data[39]~q ),
	.out_data_40(\avalon_st_adapter|data_format_adapter_0|out_data[40]~q ),
	.out_data_41(\avalon_st_adapter|data_format_adapter_0|out_data[41]~q ),
	.out_data_42(\avalon_st_adapter|data_format_adapter_0|out_data[42]~q ),
	.out_data_43(\avalon_st_adapter|data_format_adapter_0|out_data[43]~q ),
	.out_data_44(\avalon_st_adapter|data_format_adapter_0|out_data[44]~q ),
	.out_data_45(\avalon_st_adapter|data_format_adapter_0|out_data[45]~q ),
	.out_data_46(\avalon_st_adapter|data_format_adapter_0|out_data[46]~q ),
	.out_data_47(\avalon_st_adapter|data_format_adapter_0|out_data[47]~q ),
	.out_valid(\avalon_st_adapter|data_format_adapter_0|out_valid~q ),
	.avalon_streaming_source_data_0(\packet_presence_detection_0|avalon_streaming_source_data[0]~1_combout ),
	.avalon_streaming_source_data_1(\packet_presence_detection_0|avalon_streaming_source_data[1]~2_combout ),
	.avalon_streaming_source_data_2(\packet_presence_detection_0|avalon_streaming_source_data[2]~3_combout ),
	.avalon_streaming_source_data_3(\packet_presence_detection_0|avalon_streaming_source_data[3]~4_combout ),
	.avalon_streaming_source_data_4(\packet_presence_detection_0|avalon_streaming_source_data[4]~5_combout ),
	.avalon_streaming_source_data_5(\packet_presence_detection_0|avalon_streaming_source_data[5]~6_combout ),
	.avalon_streaming_source_data_6(\packet_presence_detection_0|avalon_streaming_source_data[6]~7_combout ),
	.avalon_streaming_source_data_7(\packet_presence_detection_0|avalon_streaming_source_data[7]~8_combout ),
	.avalon_streaming_source_data_8(\packet_presence_detection_0|avalon_streaming_source_data[8]~9_combout ),
	.avalon_streaming_source_data_9(\packet_presence_detection_0|avalon_streaming_source_data[9]~10_combout ),
	.avalon_streaming_source_data_10(\packet_presence_detection_0|avalon_streaming_source_data[10]~11_combout ),
	.avalon_streaming_source_data_11(\packet_presence_detection_0|avalon_streaming_source_data[11]~12_combout ),
	.avalon_streaming_source_data_12(\packet_presence_detection_0|avalon_streaming_source_data[12]~13_combout ),
	.avalon_streaming_source_data_13(\packet_presence_detection_0|avalon_streaming_source_data[13]~14_combout ),
	.avalon_streaming_source_data_14(\packet_presence_detection_0|avalon_streaming_source_data[14]~15_combout ),
	.avalon_streaming_source_data_15(\packet_presence_detection_0|avalon_streaming_source_data[15]~16_combout ),
	.avalon_streaming_source_data_16(\packet_presence_detection_0|avalon_streaming_source_data[16]~17_combout ),
	.avalon_streaming_source_data_17(\packet_presence_detection_0|avalon_streaming_source_data[17]~18_combout ),
	.avalon_streaming_source_data_18(\packet_presence_detection_0|avalon_streaming_source_data[18]~19_combout ),
	.avalon_streaming_source_data_19(\packet_presence_detection_0|avalon_streaming_source_data[19]~20_combout ),
	.avalon_streaming_source_data_20(\packet_presence_detection_0|avalon_streaming_source_data[20]~21_combout ),
	.avalon_streaming_source_data_21(\packet_presence_detection_0|avalon_streaming_source_data[21]~22_combout ),
	.avalon_streaming_source_data_22(\packet_presence_detection_0|avalon_streaming_source_data[22]~23_combout ),
	.avalon_streaming_source_data_23(\packet_presence_detection_0|avalon_streaming_source_data[23]~24_combout ),
	.delay_reg_24_3(\packet_presence_detection_0|delay_line_inst|delay_reg[3][24]~q ),
	.clk_clk(\clk_clk~input_o ));

lms_dsp_packet_presence_detection packet_presence_detection_0(
	.count_reg_0(\packet_presence_detection_0|counter_inst|count_reg[0]~q ),
	.short_sum_reg_0(\packet_presence_detection_0|running_sum_inst|short_sum_reg[0]~q ),
	.short_sum_reg_1(\packet_presence_detection_0|running_sum_inst|short_sum_reg[1]~q ),
	.short_sum_reg_2(\packet_presence_detection_0|running_sum_inst|short_sum_reg[2]~q ),
	.short_sum_reg_3(\packet_presence_detection_0|running_sum_inst|short_sum_reg[3]~q ),
	.short_sum_reg_4(\packet_presence_detection_0|running_sum_inst|short_sum_reg[4]~q ),
	.short_sum_reg_5(\packet_presence_detection_0|running_sum_inst|short_sum_reg[5]~q ),
	.short_sum_reg_6(\packet_presence_detection_0|running_sum_inst|short_sum_reg[6]~q ),
	.short_sum_reg_7(\packet_presence_detection_0|running_sum_inst|short_sum_reg[7]~q ),
	.short_sum_reg_8(\packet_presence_detection_0|running_sum_inst|short_sum_reg[8]~q ),
	.short_sum_reg_9(\packet_presence_detection_0|running_sum_inst|short_sum_reg[9]~q ),
	.short_sum_reg_10(\packet_presence_detection_0|running_sum_inst|short_sum_reg[10]~q ),
	.short_sum_reg_11(\packet_presence_detection_0|running_sum_inst|short_sum_reg[11]~q ),
	.short_sum_reg_12(\packet_presence_detection_0|running_sum_inst|short_sum_reg[12]~q ),
	.short_sum_reg_13(\packet_presence_detection_0|running_sum_inst|short_sum_reg[13]~q ),
	.short_sum_reg_14(\packet_presence_detection_0|running_sum_inst|short_sum_reg[14]~q ),
	.short_sum_reg_15(\packet_presence_detection_0|running_sum_inst|short_sum_reg[15]~q ),
	.short_sum_reg_16(\packet_presence_detection_0|running_sum_inst|short_sum_reg[16]~q ),
	.short_sum_reg_17(\packet_presence_detection_0|running_sum_inst|short_sum_reg[17]~q ),
	.count_reg_1(\packet_presence_detection_0|counter_inst|count_reg[1]~q ),
	.count_reg_2(\packet_presence_detection_0|counter_inst|count_reg[2]~q ),
	.count_reg_3(\packet_presence_detection_0|counter_inst|count_reg[3]~q ),
	.count_reg_4(\packet_presence_detection_0|counter_inst|count_reg[4]~q ),
	.count_reg_5(\packet_presence_detection_0|counter_inst|count_reg[5]~q ),
	.count_reg_6(\packet_presence_detection_0|counter_inst|count_reg[6]~q ),
	.count_reg_7(\packet_presence_detection_0|counter_inst|count_reg[7]~q ),
	.count_reg_8(\packet_presence_detection_0|counter_inst|count_reg[8]~q ),
	.count_reg_9(\packet_presence_detection_0|counter_inst|count_reg[9]~q ),
	.count_reg_10(\packet_presence_detection_0|counter_inst|count_reg[10]~q ),
	.count_reg_11(\packet_presence_detection_0|counter_inst|count_reg[11]~q ),
	.count_reg_12(\packet_presence_detection_0|counter_inst|count_reg[12]~q ),
	.count_reg_13(\packet_presence_detection_0|counter_inst|count_reg[13]~q ),
	.count_reg_14(\packet_presence_detection_0|counter_inst|count_reg[14]~q ),
	.count_reg_15(\packet_presence_detection_0|counter_inst|count_reg[15]~q ),
	.long_shift_rescale_0(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[0]~q ),
	.long_shift_rescale_1(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[1]~q ),
	.long_shift_rescale_2(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[2]~q ),
	.long_shift_rescale_3(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[3]~q ),
	.long_shift_rescale_4(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[4]~q ),
	.long_shift_rescale_5(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[5]~q ),
	.long_shift_rescale_6(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[6]~q ),
	.long_shift_rescale_7(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[7]~q ),
	.long_shift_rescale_8(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[8]~q ),
	.long_shift_rescale_9(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[9]~q ),
	.long_shift_rescale_10(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[10]~q ),
	.long_shift_rescale_11(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[11]~q ),
	.long_shift_rescale_12(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[12]~q ),
	.long_shift_rescale_13(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[13]~q ),
	.long_shift_rescale_14(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[14]~q ),
	.long_shift_rescale_15(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[15]~q ),
	.long_shift_rescale_16(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[16]~q ),
	.long_shift_rescale_17(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[17]~q ),
	.long_shift_rescale_18(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[18]~q ),
	.long_shift_rescale_19(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[19]~q ),
	.long_shift_rescale_20(\packet_presence_detection_0|running_sum_inst|long_shift_rescale[20]~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.data_out_12(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[12]~q ),
	.data_out_0(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[0]~q ),
	.data_out_11(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[11]~q ),
	.data_out_10(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[10]~q ),
	.data_out_9(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[9]~q ),
	.data_out_8(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[8]~q ),
	.data_out_7(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[7]~q ),
	.data_out_6(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[6]~q ),
	.data_out_5(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[5]~q ),
	.data_out_4(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[4]~q ),
	.data_out_3(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[3]~q ),
	.data_out_2(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[2]~q ),
	.data_out_1(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[1]~q ),
	.data_out_23(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[23]~q ),
	.data_out_22(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[22]~q ),
	.data_out_21(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[21]~q ),
	.data_out_20(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[20]~q ),
	.data_out_19(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[19]~q ),
	.data_out_18(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[18]~q ),
	.data_out_17(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[17]~q ),
	.data_out_16(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[16]~q ),
	.data_out_15(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[15]~q ),
	.data_out_14(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[14]~q ),
	.data_out_13(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[13]~q ),
	.data_valid(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_valid~q ),
	.avalon_streaming_source_data_0(\packet_presence_detection_0|avalon_streaming_source_data[0]~1_combout ),
	.avalon_streaming_source_data_1(\packet_presence_detection_0|avalon_streaming_source_data[1]~2_combout ),
	.avalon_streaming_source_data_2(\packet_presence_detection_0|avalon_streaming_source_data[2]~3_combout ),
	.avalon_streaming_source_data_3(\packet_presence_detection_0|avalon_streaming_source_data[3]~4_combout ),
	.avalon_streaming_source_data_4(\packet_presence_detection_0|avalon_streaming_source_data[4]~5_combout ),
	.avalon_streaming_source_data_5(\packet_presence_detection_0|avalon_streaming_source_data[5]~6_combout ),
	.avalon_streaming_source_data_6(\packet_presence_detection_0|avalon_streaming_source_data[6]~7_combout ),
	.avalon_streaming_source_data_7(\packet_presence_detection_0|avalon_streaming_source_data[7]~8_combout ),
	.avalon_streaming_source_data_8(\packet_presence_detection_0|avalon_streaming_source_data[8]~9_combout ),
	.avalon_streaming_source_data_9(\packet_presence_detection_0|avalon_streaming_source_data[9]~10_combout ),
	.avalon_streaming_source_data_10(\packet_presence_detection_0|avalon_streaming_source_data[10]~11_combout ),
	.avalon_streaming_source_data_11(\packet_presence_detection_0|avalon_streaming_source_data[11]~12_combout ),
	.avalon_streaming_source_data_12(\packet_presence_detection_0|avalon_streaming_source_data[12]~13_combout ),
	.avalon_streaming_source_data_13(\packet_presence_detection_0|avalon_streaming_source_data[13]~14_combout ),
	.avalon_streaming_source_data_14(\packet_presence_detection_0|avalon_streaming_source_data[14]~15_combout ),
	.avalon_streaming_source_data_15(\packet_presence_detection_0|avalon_streaming_source_data[15]~16_combout ),
	.avalon_streaming_source_data_16(\packet_presence_detection_0|avalon_streaming_source_data[16]~17_combout ),
	.avalon_streaming_source_data_17(\packet_presence_detection_0|avalon_streaming_source_data[17]~18_combout ),
	.avalon_streaming_source_data_18(\packet_presence_detection_0|avalon_streaming_source_data[18]~19_combout ),
	.avalon_streaming_source_data_19(\packet_presence_detection_0|avalon_streaming_source_data[19]~20_combout ),
	.avalon_streaming_source_data_20(\packet_presence_detection_0|avalon_streaming_source_data[20]~21_combout ),
	.avalon_streaming_source_data_21(\packet_presence_detection_0|avalon_streaming_source_data[21]~22_combout ),
	.avalon_streaming_source_data_22(\packet_presence_detection_0|avalon_streaming_source_data[22]~23_combout ),
	.avalon_streaming_source_data_23(\packet_presence_detection_0|avalon_streaming_source_data[23]~24_combout ),
	.delay_reg_24_3(\packet_presence_detection_0|delay_line_inst|delay_reg[3][24]~q ),
	.GND_port(\~GND~combout ),
	.clk_clk(\clk_clk~input_o ),
	.ppd_cfg_passthrough_len_15(\ppd_cfg_passthrough_len[15]~input_o ),
	.ppd_cfg_passthrough_len_14(\ppd_cfg_passthrough_len[14]~input_o ),
	.ppd_cfg_passthrough_len_13(\ppd_cfg_passthrough_len[13]~input_o ),
	.ppd_cfg_passthrough_len_12(\ppd_cfg_passthrough_len[12]~input_o ),
	.ppd_cfg_passthrough_len_11(\ppd_cfg_passthrough_len[11]~input_o ),
	.ppd_cfg_passthrough_len_10(\ppd_cfg_passthrough_len[10]~input_o ),
	.ppd_cfg_passthrough_len_9(\ppd_cfg_passthrough_len[9]~input_o ),
	.ppd_cfg_passthrough_len_8(\ppd_cfg_passthrough_len[8]~input_o ),
	.ppd_cfg_passthrough_len_7(\ppd_cfg_passthrough_len[7]~input_o ),
	.ppd_cfg_passthrough_len_6(\ppd_cfg_passthrough_len[6]~input_o ),
	.ppd_cfg_passthrough_len_5(\ppd_cfg_passthrough_len[5]~input_o ),
	.ppd_cfg_passthrough_len_4(\ppd_cfg_passthrough_len[4]~input_o ),
	.ppd_cfg_passthrough_len_3(\ppd_cfg_passthrough_len[3]~input_o ),
	.ppd_cfg_passthrough_len_2(\ppd_cfg_passthrough_len[2]~input_o ),
	.ppd_cfg_passthrough_len_1(\ppd_cfg_passthrough_len[1]~input_o ),
	.ppd_cfg_passthrough_len_0(\ppd_cfg_passthrough_len[0]~input_o ),
	.ppd_cfg_clear_rs(\ppd_cfg_clear_rs~input_o ),
	.ppd_cfg_threshold_0(\ppd_cfg_threshold[0]~input_o ),
	.ppd_cfg_threshold_1(\ppd_cfg_threshold[1]~input_o ),
	.ppd_cfg_threshold_2(\ppd_cfg_threshold[2]~input_o ),
	.ppd_cfg_threshold_3(\ppd_cfg_threshold[3]~input_o ),
	.ppd_cfg_threshold_4(\ppd_cfg_threshold[4]~input_o ),
	.ppd_cfg_threshold_5(\ppd_cfg_threshold[5]~input_o ),
	.ppd_cfg_threshold_6(\ppd_cfg_threshold[6]~input_o ),
	.ppd_cfg_threshold_7(\ppd_cfg_threshold[7]~input_o ),
	.ppd_cfg_enable(\ppd_cfg_enable~input_o ));

lms_dsp_lms_dsp_fir_compiler_ii_0 fir_compiler_ii_0(
	.reset_n(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.data_out_12(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[12]~q ),
	.data_out_0(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[0]~q ),
	.data_out_11(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[11]~q ),
	.data_out_10(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[10]~q ),
	.data_out_9(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[9]~q ),
	.data_out_8(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[8]~q ),
	.data_out_7(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[7]~q ),
	.data_out_6(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[6]~q ),
	.data_out_5(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[5]~q ),
	.data_out_4(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[4]~q ),
	.data_out_3(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[3]~q ),
	.data_out_2(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[2]~q ),
	.data_out_1(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[1]~q ),
	.data_out_23(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[23]~q ),
	.data_out_22(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[22]~q ),
	.data_out_21(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[21]~q ),
	.data_out_20(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[20]~q ),
	.data_out_19(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[19]~q ),
	.data_out_18(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[18]~q ),
	.data_out_17(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[17]~q ),
	.data_out_16(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[16]~q ),
	.data_out_15(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[15]~q ),
	.data_out_14(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[14]~q ),
	.data_out_13(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_out[13]~q ),
	.data_valid(\fir_compiler_ii_0|lms_dsp_fir_compiler_ii_0_ast_inst|source|data_valid~q ),
	.out_valid(\avalon_st_adapter_001|data_format_adapter_0|out_valid~q ),
	.out_data_21(\avalon_st_adapter_001|data_format_adapter_0|out_data[21]~q ),
	.out_data_20(\avalon_st_adapter_001|data_format_adapter_0|out_data[20]~q ),
	.out_data_19(\avalon_st_adapter_001|data_format_adapter_0|out_data[19]~q ),
	.out_data_18(\avalon_st_adapter_001|data_format_adapter_0|out_data[18]~q ),
	.out_data_17(\avalon_st_adapter_001|data_format_adapter_0|out_data[17]~q ),
	.out_data_16(\avalon_st_adapter_001|data_format_adapter_0|out_data[16]~q ),
	.out_data_15(\avalon_st_adapter_001|data_format_adapter_0|out_data[15]~q ),
	.out_data_14(\avalon_st_adapter_001|data_format_adapter_0|out_data[14]~q ),
	.out_data_12(\avalon_st_adapter_001|data_format_adapter_0|out_data[12]~q ),
	.out_data_13(\avalon_st_adapter_001|data_format_adapter_0|out_data[13]~q ),
	.out_data_9(\avalon_st_adapter_001|data_format_adapter_0|out_data[9]~q ),
	.out_data_8(\avalon_st_adapter_001|data_format_adapter_0|out_data[8]~q ),
	.out_data_7(\avalon_st_adapter_001|data_format_adapter_0|out_data[7]~q ),
	.out_data_6(\avalon_st_adapter_001|data_format_adapter_0|out_data[6]~q ),
	.out_data_5(\avalon_st_adapter_001|data_format_adapter_0|out_data[5]~q ),
	.out_data_4(\avalon_st_adapter_001|data_format_adapter_0|out_data[4]~q ),
	.out_data_3(\avalon_st_adapter_001|data_format_adapter_0|out_data[3]~q ),
	.out_data_2(\avalon_st_adapter_001|data_format_adapter_0|out_data[2]~q ),
	.out_data_0(\avalon_st_adapter_001|data_format_adapter_0|out_data[0]~q ),
	.out_data_1(\avalon_st_adapter_001|data_format_adapter_0|out_data[1]~q ),
	.out_data_11(\avalon_st_adapter_001|data_format_adapter_0|out_data[11]~q ),
	.out_data_10(\avalon_st_adapter_001|data_format_adapter_0|out_data[10]~q ),
	.out_data_23(\avalon_st_adapter_001|data_format_adapter_0|out_data[23]~q ),
	.out_data_22(\avalon_st_adapter_001|data_format_adapter_0|out_data[22]~q ),
	.clk(\clk_clk~input_o ));

lms_dsp_fifo2avs fifo2avs_0(
	.reset_sink_reset(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.valid_reg1(\fifo2avs_0|valid_reg~q ),
	.data_reg_21(\fifo2avs_0|data_reg[21]~q ),
	.data_reg_45(\fifo2avs_0|data_reg[45]~q ),
	.data_reg_20(\fifo2avs_0|data_reg[20]~q ),
	.data_reg_44(\fifo2avs_0|data_reg[44]~q ),
	.data_reg_19(\fifo2avs_0|data_reg[19]~q ),
	.data_reg_43(\fifo2avs_0|data_reg[43]~q ),
	.data_reg_18(\fifo2avs_0|data_reg[18]~q ),
	.data_reg_42(\fifo2avs_0|data_reg[42]~q ),
	.data_reg_17(\fifo2avs_0|data_reg[17]~q ),
	.data_reg_41(\fifo2avs_0|data_reg[41]~q ),
	.data_reg_16(\fifo2avs_0|data_reg[16]~q ),
	.data_reg_40(\fifo2avs_0|data_reg[40]~q ),
	.data_reg_15(\fifo2avs_0|data_reg[15]~q ),
	.data_reg_39(\fifo2avs_0|data_reg[39]~q ),
	.data_reg_14(\fifo2avs_0|data_reg[14]~q ),
	.data_reg_38(\fifo2avs_0|data_reg[38]~q ),
	.data_reg_12(\fifo2avs_0|data_reg[12]~q ),
	.data_reg_36(\fifo2avs_0|data_reg[36]~q ),
	.data_reg_13(\fifo2avs_0|data_reg[13]~q ),
	.data_reg_37(\fifo2avs_0|data_reg[37]~q ),
	.data_reg_9(\fifo2avs_0|data_reg[9]~q ),
	.data_reg_33(\fifo2avs_0|data_reg[33]~q ),
	.data_reg_8(\fifo2avs_0|data_reg[8]~q ),
	.data_reg_32(\fifo2avs_0|data_reg[32]~q ),
	.data_reg_7(\fifo2avs_0|data_reg[7]~q ),
	.data_reg_31(\fifo2avs_0|data_reg[31]~q ),
	.data_reg_6(\fifo2avs_0|data_reg[6]~q ),
	.data_reg_30(\fifo2avs_0|data_reg[30]~q ),
	.data_reg_5(\fifo2avs_0|data_reg[5]~q ),
	.data_reg_29(\fifo2avs_0|data_reg[29]~q ),
	.data_reg_4(\fifo2avs_0|data_reg[4]~q ),
	.data_reg_28(\fifo2avs_0|data_reg[28]~q ),
	.data_reg_3(\fifo2avs_0|data_reg[3]~q ),
	.data_reg_27(\fifo2avs_0|data_reg[27]~q ),
	.data_reg_2(\fifo2avs_0|data_reg[2]~q ),
	.data_reg_26(\fifo2avs_0|data_reg[26]~q ),
	.data_reg_0(\fifo2avs_0|data_reg[0]~q ),
	.data_reg_24(\fifo2avs_0|data_reg[24]~q ),
	.data_reg_1(\fifo2avs_0|data_reg[1]~q ),
	.data_reg_25(\fifo2avs_0|data_reg[25]~q ),
	.data_reg_11(\fifo2avs_0|data_reg[11]~q ),
	.data_reg_35(\fifo2avs_0|data_reg[35]~q ),
	.data_reg_10(\fifo2avs_0|data_reg[10]~q ),
	.data_reg_34(\fifo2avs_0|data_reg[34]~q ),
	.data_reg_23(\fifo2avs_0|data_reg[23]~q ),
	.data_reg_47(\fifo2avs_0|data_reg[47]~q ),
	.data_reg_22(\fifo2avs_0|data_reg[22]~q ),
	.data_reg_46(\fifo2avs_0|data_reg[46]~q ),
	.clock_sink_clk(\clk_clk~input_o ),
	.fifo_wrreq(\fifo_in_wrreq~input_o ),
	.fifo_wdata({\fifo_in_wdata[47]~input_o ,\fifo_in_wdata[46]~input_o ,\fifo_in_wdata[45]~input_o ,\fifo_in_wdata[44]~input_o ,\fifo_in_wdata[43]~input_o ,\fifo_in_wdata[42]~input_o ,\fifo_in_wdata[41]~input_o ,\fifo_in_wdata[40]~input_o ,\fifo_in_wdata[39]~input_o ,
\fifo_in_wdata[38]~input_o ,\fifo_in_wdata[37]~input_o ,\fifo_in_wdata[36]~input_o ,\fifo_in_wdata[35]~input_o ,\fifo_in_wdata[34]~input_o ,\fifo_in_wdata[33]~input_o ,\fifo_in_wdata[32]~input_o ,\fifo_in_wdata[31]~input_o ,\fifo_in_wdata[30]~input_o ,
\fifo_in_wdata[29]~input_o ,\fifo_in_wdata[28]~input_o ,\fifo_in_wdata[27]~input_o ,\fifo_in_wdata[26]~input_o ,\fifo_in_wdata[25]~input_o ,\fifo_in_wdata[24]~input_o ,\fifo_in_wdata[23]~input_o ,\fifo_in_wdata[22]~input_o ,\fifo_in_wdata[21]~input_o ,
\fifo_in_wdata[20]~input_o ,\fifo_in_wdata[19]~input_o ,\fifo_in_wdata[18]~input_o ,\fifo_in_wdata[17]~input_o ,\fifo_in_wdata[16]~input_o ,\fifo_in_wdata[15]~input_o ,\fifo_in_wdata[14]~input_o ,\fifo_in_wdata[13]~input_o ,\fifo_in_wdata[12]~input_o ,
\fifo_in_wdata[11]~input_o ,\fifo_in_wdata[10]~input_o ,\fifo_in_wdata[9]~input_o ,\fifo_in_wdata[8]~input_o ,\fifo_in_wdata[7]~input_o ,\fifo_in_wdata[6]~input_o ,\fifo_in_wdata[5]~input_o ,\fifo_in_wdata[4]~input_o ,\fifo_in_wdata[3]~input_o ,
\fifo_in_wdata[2]~input_o ,\fifo_in_wdata[1]~input_o ,\fifo_in_wdata[0]~input_o }));

lms_dsp_avs2fifo avs2fifo_0(
	.wrdata_reg_0(\avs2fifo_0|wrdata_reg[0]~q ),
	.wrdata_reg_1(\avs2fifo_0|wrdata_reg[1]~q ),
	.wrdata_reg_2(\avs2fifo_0|wrdata_reg[2]~q ),
	.wrdata_reg_3(\avs2fifo_0|wrdata_reg[3]~q ),
	.wrdata_reg_4(\avs2fifo_0|wrdata_reg[4]~q ),
	.wrdata_reg_5(\avs2fifo_0|wrdata_reg[5]~q ),
	.wrdata_reg_6(\avs2fifo_0|wrdata_reg[6]~q ),
	.wrdata_reg_7(\avs2fifo_0|wrdata_reg[7]~q ),
	.wrdata_reg_8(\avs2fifo_0|wrdata_reg[8]~q ),
	.wrdata_reg_9(\avs2fifo_0|wrdata_reg[9]~q ),
	.wrdata_reg_10(\avs2fifo_0|wrdata_reg[10]~q ),
	.wrdata_reg_11(\avs2fifo_0|wrdata_reg[11]~q ),
	.wrdata_reg_12(\avs2fifo_0|wrdata_reg[12]~q ),
	.wrdata_reg_13(\avs2fifo_0|wrdata_reg[13]~q ),
	.wrdata_reg_14(\avs2fifo_0|wrdata_reg[14]~q ),
	.wrdata_reg_15(\avs2fifo_0|wrdata_reg[15]~q ),
	.wrdata_reg_16(\avs2fifo_0|wrdata_reg[16]~q ),
	.wrdata_reg_17(\avs2fifo_0|wrdata_reg[17]~q ),
	.wrdata_reg_18(\avs2fifo_0|wrdata_reg[18]~q ),
	.wrdata_reg_19(\avs2fifo_0|wrdata_reg[19]~q ),
	.wrdata_reg_20(\avs2fifo_0|wrdata_reg[20]~q ),
	.wrdata_reg_21(\avs2fifo_0|wrdata_reg[21]~q ),
	.wrdata_reg_22(\avs2fifo_0|wrdata_reg[22]~q ),
	.wrdata_reg_23(\avs2fifo_0|wrdata_reg[23]~q ),
	.wrdata_reg_24(\avs2fifo_0|wrdata_reg[24]~q ),
	.wrdata_reg_25(\avs2fifo_0|wrdata_reg[25]~q ),
	.wrdata_reg_26(\avs2fifo_0|wrdata_reg[26]~q ),
	.wrdata_reg_27(\avs2fifo_0|wrdata_reg[27]~q ),
	.wrdata_reg_28(\avs2fifo_0|wrdata_reg[28]~q ),
	.wrdata_reg_29(\avs2fifo_0|wrdata_reg[29]~q ),
	.wrdata_reg_30(\avs2fifo_0|wrdata_reg[30]~q ),
	.wrdata_reg_31(\avs2fifo_0|wrdata_reg[31]~q ),
	.wrdata_reg_32(\avs2fifo_0|wrdata_reg[32]~q ),
	.wrdata_reg_33(\avs2fifo_0|wrdata_reg[33]~q ),
	.wrdata_reg_34(\avs2fifo_0|wrdata_reg[34]~q ),
	.wrdata_reg_35(\avs2fifo_0|wrdata_reg[35]~q ),
	.wrdata_reg_36(\avs2fifo_0|wrdata_reg[36]~q ),
	.wrdata_reg_37(\avs2fifo_0|wrdata_reg[37]~q ),
	.wrdata_reg_38(\avs2fifo_0|wrdata_reg[38]~q ),
	.wrdata_reg_39(\avs2fifo_0|wrdata_reg[39]~q ),
	.wrdata_reg_40(\avs2fifo_0|wrdata_reg[40]~q ),
	.wrdata_reg_41(\avs2fifo_0|wrdata_reg[41]~q ),
	.wrdata_reg_42(\avs2fifo_0|wrdata_reg[42]~q ),
	.wrdata_reg_43(\avs2fifo_0|wrdata_reg[43]~q ),
	.wrdata_reg_44(\avs2fifo_0|wrdata_reg[44]~q ),
	.wrdata_reg_45(\avs2fifo_0|wrdata_reg[45]~q ),
	.wrdata_reg_46(\avs2fifo_0|wrdata_reg[46]~q ),
	.wrdata_reg_47(\avs2fifo_0|wrdata_reg[47]~q ),
	.wrreq_reg1(\avs2fifo_0|wrreq_reg~q ),
	.avalon_streaming_sink_data({\avalon_st_adapter|data_format_adapter_0|out_data[47]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[46]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[45]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[44]~q ,
\avalon_st_adapter|data_format_adapter_0|out_data[43]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[42]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[41]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[40]~q ,
\avalon_st_adapter|data_format_adapter_0|out_data[39]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[38]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[37]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[36]~q ,
\avalon_st_adapter|data_format_adapter_0|out_data[35]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[34]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[33]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[32]~q ,
\avalon_st_adapter|data_format_adapter_0|out_data[31]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[30]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[29]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[28]~q ,
\avalon_st_adapter|data_format_adapter_0|out_data[27]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[26]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[25]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[24]~q ,
\avalon_st_adapter|data_format_adapter_0|out_data[23]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[22]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[21]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[20]~q ,
\avalon_st_adapter|data_format_adapter_0|out_data[19]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[18]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[17]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[16]~q ,
\avalon_st_adapter|data_format_adapter_0|out_data[15]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[14]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[13]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[12]~q ,
\avalon_st_adapter|data_format_adapter_0|out_data[11]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[10]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[9]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[8]~q ,
\avalon_st_adapter|data_format_adapter_0|out_data[7]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[6]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[5]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[4]~q ,
\avalon_st_adapter|data_format_adapter_0|out_data[3]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[2]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[1]~q ,\avalon_st_adapter|data_format_adapter_0|out_data[0]~q }),
	.reset_sink_reset(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.avalon_streaming_sink_valid(\avalon_st_adapter|data_format_adapter_0|out_valid~q ),
	.clock_sink_clk(\clk_clk~input_o ));

fiftyfivenm_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~GND~combout ),
	.cout());
defparam \~GND .lut_mask = 16'h0000;
defparam \~GND .sum_lutc_input = "datac";

assign \clk_clk~input_o  = clk_clk;

assign \ppd_cfg_passthrough_len[15]~input_o  = ppd_cfg_passthrough_len[15];

assign \ppd_cfg_passthrough_len[14]~input_o  = ppd_cfg_passthrough_len[14];

assign \ppd_cfg_passthrough_len[13]~input_o  = ppd_cfg_passthrough_len[13];

assign \ppd_cfg_passthrough_len[12]~input_o  = ppd_cfg_passthrough_len[12];

assign \ppd_cfg_passthrough_len[11]~input_o  = ppd_cfg_passthrough_len[11];

assign \ppd_cfg_passthrough_len[10]~input_o  = ppd_cfg_passthrough_len[10];

assign \ppd_cfg_passthrough_len[9]~input_o  = ppd_cfg_passthrough_len[9];

assign \ppd_cfg_passthrough_len[8]~input_o  = ppd_cfg_passthrough_len[8];

assign \ppd_cfg_passthrough_len[7]~input_o  = ppd_cfg_passthrough_len[7];

assign \ppd_cfg_passthrough_len[6]~input_o  = ppd_cfg_passthrough_len[6];

assign \ppd_cfg_passthrough_len[5]~input_o  = ppd_cfg_passthrough_len[5];

assign \ppd_cfg_passthrough_len[4]~input_o  = ppd_cfg_passthrough_len[4];

assign \ppd_cfg_passthrough_len[3]~input_o  = ppd_cfg_passthrough_len[3];

assign \ppd_cfg_passthrough_len[2]~input_o  = ppd_cfg_passthrough_len[2];

assign \ppd_cfg_passthrough_len[1]~input_o  = ppd_cfg_passthrough_len[1];

assign \ppd_cfg_passthrough_len[0]~input_o  = ppd_cfg_passthrough_len[0];

assign \ppd_cfg_clear_rs~input_o  = ppd_cfg_clear_rs;

assign \reset_reset_n~input_o  = reset_reset_n;

assign \ppd_cfg_threshold[0]~input_o  = ppd_cfg_threshold[0];

assign \ppd_cfg_threshold[1]~input_o  = ppd_cfg_threshold[1];

assign \ppd_cfg_threshold[2]~input_o  = ppd_cfg_threshold[2];

assign \ppd_cfg_threshold[3]~input_o  = ppd_cfg_threshold[3];

assign \ppd_cfg_threshold[4]~input_o  = ppd_cfg_threshold[4];

assign \ppd_cfg_threshold[5]~input_o  = ppd_cfg_threshold[5];

assign \ppd_cfg_threshold[6]~input_o  = ppd_cfg_threshold[6];

assign \ppd_cfg_threshold[7]~input_o  = ppd_cfg_threshold[7];

assign \ppd_cfg_enable~input_o  = ppd_cfg_enable;

assign \fifo_in_wrreq~input_o  = fifo_in_wrreq;

assign \fifo_in_wdata[21]~input_o  = fifo_in_wdata[21];

assign \fifo_in_wdata[45]~input_o  = fifo_in_wdata[45];

assign \fifo_in_wdata[20]~input_o  = fifo_in_wdata[20];

assign \fifo_in_wdata[44]~input_o  = fifo_in_wdata[44];

assign \fifo_in_wdata[19]~input_o  = fifo_in_wdata[19];

assign \fifo_in_wdata[43]~input_o  = fifo_in_wdata[43];

assign \fifo_in_wdata[18]~input_o  = fifo_in_wdata[18];

assign \fifo_in_wdata[42]~input_o  = fifo_in_wdata[42];

assign \fifo_in_wdata[17]~input_o  = fifo_in_wdata[17];

assign \fifo_in_wdata[41]~input_o  = fifo_in_wdata[41];

assign \fifo_in_wdata[16]~input_o  = fifo_in_wdata[16];

assign \fifo_in_wdata[40]~input_o  = fifo_in_wdata[40];

assign \fifo_in_wdata[15]~input_o  = fifo_in_wdata[15];

assign \fifo_in_wdata[39]~input_o  = fifo_in_wdata[39];

assign \fifo_in_wdata[14]~input_o  = fifo_in_wdata[14];

assign \fifo_in_wdata[38]~input_o  = fifo_in_wdata[38];

assign \fifo_in_wdata[12]~input_o  = fifo_in_wdata[12];

assign \fifo_in_wdata[36]~input_o  = fifo_in_wdata[36];

assign \fifo_in_wdata[13]~input_o  = fifo_in_wdata[13];

assign \fifo_in_wdata[37]~input_o  = fifo_in_wdata[37];

assign \fifo_in_wdata[9]~input_o  = fifo_in_wdata[9];

assign \fifo_in_wdata[33]~input_o  = fifo_in_wdata[33];

assign \fifo_in_wdata[8]~input_o  = fifo_in_wdata[8];

assign \fifo_in_wdata[32]~input_o  = fifo_in_wdata[32];

assign \fifo_in_wdata[7]~input_o  = fifo_in_wdata[7];

assign \fifo_in_wdata[31]~input_o  = fifo_in_wdata[31];

assign \fifo_in_wdata[6]~input_o  = fifo_in_wdata[6];

assign \fifo_in_wdata[30]~input_o  = fifo_in_wdata[30];

assign \fifo_in_wdata[5]~input_o  = fifo_in_wdata[5];

assign \fifo_in_wdata[29]~input_o  = fifo_in_wdata[29];

assign \fifo_in_wdata[4]~input_o  = fifo_in_wdata[4];

assign \fifo_in_wdata[28]~input_o  = fifo_in_wdata[28];

assign \fifo_in_wdata[3]~input_o  = fifo_in_wdata[3];

assign \fifo_in_wdata[27]~input_o  = fifo_in_wdata[27];

assign \fifo_in_wdata[2]~input_o  = fifo_in_wdata[2];

assign \fifo_in_wdata[26]~input_o  = fifo_in_wdata[26];

assign \fifo_in_wdata[0]~input_o  = fifo_in_wdata[0];

assign \fifo_in_wdata[24]~input_o  = fifo_in_wdata[24];

assign \fifo_in_wdata[1]~input_o  = fifo_in_wdata[1];

assign \fifo_in_wdata[25]~input_o  = fifo_in_wdata[25];

assign \fifo_in_wdata[11]~input_o  = fifo_in_wdata[11];

assign \fifo_in_wdata[35]~input_o  = fifo_in_wdata[35];

assign \fifo_in_wdata[10]~input_o  = fifo_in_wdata[10];

assign \fifo_in_wdata[34]~input_o  = fifo_in_wdata[34];

assign \fifo_in_wdata[23]~input_o  = fifo_in_wdata[23];

assign \fifo_in_wdata[47]~input_o  = fifo_in_wdata[47];

assign \fifo_in_wdata[22]~input_o  = fifo_in_wdata[22];

assign \fifo_in_wdata[46]~input_o  = fifo_in_wdata[46];

assign fifo_out_wrdata[0] = \avs2fifo_0|wrdata_reg[0]~q ;

assign fifo_out_wrdata[1] = \avs2fifo_0|wrdata_reg[1]~q ;

assign fifo_out_wrdata[2] = \avs2fifo_0|wrdata_reg[2]~q ;

assign fifo_out_wrdata[3] = \avs2fifo_0|wrdata_reg[3]~q ;

assign fifo_out_wrdata[4] = \avs2fifo_0|wrdata_reg[4]~q ;

assign fifo_out_wrdata[5] = \avs2fifo_0|wrdata_reg[5]~q ;

assign fifo_out_wrdata[6] = \avs2fifo_0|wrdata_reg[6]~q ;

assign fifo_out_wrdata[7] = \avs2fifo_0|wrdata_reg[7]~q ;

assign fifo_out_wrdata[8] = \avs2fifo_0|wrdata_reg[8]~q ;

assign fifo_out_wrdata[9] = \avs2fifo_0|wrdata_reg[9]~q ;

assign fifo_out_wrdata[10] = \avs2fifo_0|wrdata_reg[10]~q ;

assign fifo_out_wrdata[11] = \avs2fifo_0|wrdata_reg[11]~q ;

assign fifo_out_wrdata[12] = \avs2fifo_0|wrdata_reg[12]~q ;

assign fifo_out_wrdata[13] = \avs2fifo_0|wrdata_reg[13]~q ;

assign fifo_out_wrdata[14] = \avs2fifo_0|wrdata_reg[14]~q ;

assign fifo_out_wrdata[15] = \avs2fifo_0|wrdata_reg[15]~q ;

assign fifo_out_wrdata[16] = \avs2fifo_0|wrdata_reg[16]~q ;

assign fifo_out_wrdata[17] = \avs2fifo_0|wrdata_reg[17]~q ;

assign fifo_out_wrdata[18] = \avs2fifo_0|wrdata_reg[18]~q ;

assign fifo_out_wrdata[19] = \avs2fifo_0|wrdata_reg[19]~q ;

assign fifo_out_wrdata[20] = \avs2fifo_0|wrdata_reg[20]~q ;

assign fifo_out_wrdata[21] = \avs2fifo_0|wrdata_reg[21]~q ;

assign fifo_out_wrdata[22] = \avs2fifo_0|wrdata_reg[22]~q ;

assign fifo_out_wrdata[23] = \avs2fifo_0|wrdata_reg[23]~q ;

assign fifo_out_wrdata[24] = \avs2fifo_0|wrdata_reg[24]~q ;

assign fifo_out_wrdata[25] = \avs2fifo_0|wrdata_reg[25]~q ;

assign fifo_out_wrdata[26] = \avs2fifo_0|wrdata_reg[26]~q ;

assign fifo_out_wrdata[27] = \avs2fifo_0|wrdata_reg[27]~q ;

assign fifo_out_wrdata[28] = \avs2fifo_0|wrdata_reg[28]~q ;

assign fifo_out_wrdata[29] = \avs2fifo_0|wrdata_reg[29]~q ;

assign fifo_out_wrdata[30] = \avs2fifo_0|wrdata_reg[30]~q ;

assign fifo_out_wrdata[31] = \avs2fifo_0|wrdata_reg[31]~q ;

assign fifo_out_wrdata[32] = \avs2fifo_0|wrdata_reg[32]~q ;

assign fifo_out_wrdata[33] = \avs2fifo_0|wrdata_reg[33]~q ;

assign fifo_out_wrdata[34] = \avs2fifo_0|wrdata_reg[34]~q ;

assign fifo_out_wrdata[35] = \avs2fifo_0|wrdata_reg[35]~q ;

assign fifo_out_wrdata[36] = \avs2fifo_0|wrdata_reg[36]~q ;

assign fifo_out_wrdata[37] = \avs2fifo_0|wrdata_reg[37]~q ;

assign fifo_out_wrdata[38] = \avs2fifo_0|wrdata_reg[38]~q ;

assign fifo_out_wrdata[39] = \avs2fifo_0|wrdata_reg[39]~q ;

assign fifo_out_wrdata[40] = \avs2fifo_0|wrdata_reg[40]~q ;

assign fifo_out_wrdata[41] = \avs2fifo_0|wrdata_reg[41]~q ;

assign fifo_out_wrdata[42] = \avs2fifo_0|wrdata_reg[42]~q ;

assign fifo_out_wrdata[43] = \avs2fifo_0|wrdata_reg[43]~q ;

assign fifo_out_wrdata[44] = \avs2fifo_0|wrdata_reg[44]~q ;

assign fifo_out_wrdata[45] = \avs2fifo_0|wrdata_reg[45]~q ;

assign fifo_out_wrdata[46] = \avs2fifo_0|wrdata_reg[46]~q ;

assign fifo_out_wrdata[47] = \avs2fifo_0|wrdata_reg[47]~q ;

assign fifo_out_wrreq = \avs2fifo_0|wrreq_reg~q ;

assign ppd_debug_count[0] = \packet_presence_detection_0|counter_inst|count_reg[0]~q ;

assign ppd_debug_count[1] = \packet_presence_detection_0|counter_inst|count_reg[1]~q ;

assign ppd_debug_count[2] = \packet_presence_detection_0|counter_inst|count_reg[2]~q ;

assign ppd_debug_count[3] = \packet_presence_detection_0|counter_inst|count_reg[3]~q ;

assign ppd_debug_count[4] = \packet_presence_detection_0|counter_inst|count_reg[4]~q ;

assign ppd_debug_count[5] = \packet_presence_detection_0|counter_inst|count_reg[5]~q ;

assign ppd_debug_count[6] = \packet_presence_detection_0|counter_inst|count_reg[6]~q ;

assign ppd_debug_count[7] = \packet_presence_detection_0|counter_inst|count_reg[7]~q ;

assign ppd_debug_count[8] = \packet_presence_detection_0|counter_inst|count_reg[8]~q ;

assign ppd_debug_count[9] = \packet_presence_detection_0|counter_inst|count_reg[9]~q ;

assign ppd_debug_count[10] = \packet_presence_detection_0|counter_inst|count_reg[10]~q ;

assign ppd_debug_count[11] = \packet_presence_detection_0|counter_inst|count_reg[11]~q ;

assign ppd_debug_count[12] = \packet_presence_detection_0|counter_inst|count_reg[12]~q ;

assign ppd_debug_count[13] = \packet_presence_detection_0|counter_inst|count_reg[13]~q ;

assign ppd_debug_count[14] = \packet_presence_detection_0|counter_inst|count_reg[14]~q ;

assign ppd_debug_count[15] = \packet_presence_detection_0|counter_inst|count_reg[15]~q ;

assign ppd_debug_count[16] = gnd;

assign ppd_debug_count[17] = gnd;

assign ppd_debug_count[18] = gnd;

assign ppd_debug_count[19] = gnd;

assign ppd_debug_count[20] = gnd;

assign ppd_debug_count[21] = gnd;

assign ppd_debug_count[22] = gnd;

assign ppd_debug_count[23] = gnd;

assign ppd_debug_count[24] = gnd;

assign ppd_debug_count[25] = gnd;

assign ppd_debug_count[26] = gnd;

assign ppd_debug_count[27] = gnd;

assign ppd_debug_count[28] = gnd;

assign ppd_debug_count[29] = gnd;

assign ppd_debug_count[30] = gnd;

assign ppd_debug_count[31] = gnd;

assign ppd_debug_long_sum[0] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[0]~q ;

assign ppd_debug_long_sum[1] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[1]~q ;

assign ppd_debug_long_sum[2] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[2]~q ;

assign ppd_debug_long_sum[3] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[3]~q ;

assign ppd_debug_long_sum[4] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[4]~q ;

assign ppd_debug_long_sum[5] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[5]~q ;

assign ppd_debug_long_sum[6] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[6]~q ;

assign ppd_debug_long_sum[7] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[7]~q ;

assign ppd_debug_long_sum[8] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[8]~q ;

assign ppd_debug_long_sum[9] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[9]~q ;

assign ppd_debug_long_sum[10] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[10]~q ;

assign ppd_debug_long_sum[11] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[11]~q ;

assign ppd_debug_long_sum[12] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[12]~q ;

assign ppd_debug_long_sum[13] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[13]~q ;

assign ppd_debug_long_sum[14] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[14]~q ;

assign ppd_debug_long_sum[15] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[15]~q ;

assign ppd_debug_long_sum[16] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[16]~q ;

assign ppd_debug_long_sum[17] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[17]~q ;

assign ppd_debug_long_sum[18] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[18]~q ;

assign ppd_debug_long_sum[19] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[19]~q ;

assign ppd_debug_long_sum[20] = \packet_presence_detection_0|running_sum_inst|long_shift_rescale[20]~q ;

assign ppd_debug_long_sum[21] = gnd;

assign ppd_debug_long_sum[22] = gnd;

assign ppd_debug_long_sum[23] = gnd;

assign ppd_debug_long_sum[24] = gnd;

assign ppd_debug_long_sum[25] = gnd;

assign ppd_debug_long_sum[26] = gnd;

assign ppd_debug_long_sum[27] = gnd;

assign ppd_debug_long_sum[28] = gnd;

assign ppd_debug_long_sum[29] = gnd;

assign ppd_debug_long_sum[30] = gnd;

assign ppd_debug_long_sum[31] = gnd;

assign ppd_debug_short_sum[0] = \packet_presence_detection_0|running_sum_inst|short_sum_reg[0]~q ;

assign ppd_debug_short_sum[1] = \packet_presence_detection_0|running_sum_inst|short_sum_reg[1]~q ;

assign ppd_debug_short_sum[2] = \packet_presence_detection_0|running_sum_inst|short_sum_reg[2]~q ;

assign ppd_debug_short_sum[3] = \packet_presence_detection_0|running_sum_inst|short_sum_reg[3]~q ;

assign ppd_debug_short_sum[4] = \packet_presence_detection_0|running_sum_inst|short_sum_reg[4]~q ;

assign ppd_debug_short_sum[5] = \packet_presence_detection_0|running_sum_inst|short_sum_reg[5]~q ;

assign ppd_debug_short_sum[6] = \packet_presence_detection_0|running_sum_inst|short_sum_reg[6]~q ;

assign ppd_debug_short_sum[7] = \packet_presence_detection_0|running_sum_inst|short_sum_reg[7]~q ;

assign ppd_debug_short_sum[8] = \packet_presence_detection_0|running_sum_inst|short_sum_reg[8]~q ;

assign ppd_debug_short_sum[9] = \packet_presence_detection_0|running_sum_inst|short_sum_reg[9]~q ;

assign ppd_debug_short_sum[10] = \packet_presence_detection_0|running_sum_inst|short_sum_reg[10]~q ;

assign ppd_debug_short_sum[11] = \packet_presence_detection_0|running_sum_inst|short_sum_reg[11]~q ;

assign ppd_debug_short_sum[12] = \packet_presence_detection_0|running_sum_inst|short_sum_reg[12]~q ;

assign ppd_debug_short_sum[13] = \packet_presence_detection_0|running_sum_inst|short_sum_reg[13]~q ;

assign ppd_debug_short_sum[14] = \packet_presence_detection_0|running_sum_inst|short_sum_reg[14]~q ;

assign ppd_debug_short_sum[15] = \packet_presence_detection_0|running_sum_inst|short_sum_reg[15]~q ;

assign ppd_debug_short_sum[16] = \packet_presence_detection_0|running_sum_inst|short_sum_reg[16]~q ;

assign ppd_debug_short_sum[17] = \packet_presence_detection_0|running_sum_inst|short_sum_reg[17]~q ;

assign ppd_debug_short_sum[18] = gnd;

assign ppd_debug_short_sum[19] = gnd;

assign ppd_debug_short_sum[20] = gnd;

assign ppd_debug_short_sum[21] = gnd;

assign ppd_debug_short_sum[22] = gnd;

assign ppd_debug_short_sum[23] = gnd;

assign ppd_debug_short_sum[24] = gnd;

assign ppd_debug_short_sum[25] = gnd;

assign ppd_debug_short_sum[26] = gnd;

assign ppd_debug_short_sum[27] = gnd;

assign ppd_debug_short_sum[28] = gnd;

assign ppd_debug_short_sum[29] = gnd;

assign ppd_debug_short_sum[30] = gnd;

assign ppd_debug_short_sum[31] = gnd;

endmodule

module lms_dsp_altera_reset_controller (
	altera_reset_synchronizer_int_chain_out,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
output 	altera_reset_synchronizer_int_chain_out;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



lms_dsp_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk),
	.reset_reset_n(reset_reset_n));

endmodule

module lms_dsp_altera_reset_synchronizer_1 (
	altera_reset_synchronizer_int_chain_out1,
	clk,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module lms_dsp_avs2fifo (
	wrdata_reg_0,
	wrdata_reg_1,
	wrdata_reg_2,
	wrdata_reg_3,
	wrdata_reg_4,
	wrdata_reg_5,
	wrdata_reg_6,
	wrdata_reg_7,
	wrdata_reg_8,
	wrdata_reg_9,
	wrdata_reg_10,
	wrdata_reg_11,
	wrdata_reg_12,
	wrdata_reg_13,
	wrdata_reg_14,
	wrdata_reg_15,
	wrdata_reg_16,
	wrdata_reg_17,
	wrdata_reg_18,
	wrdata_reg_19,
	wrdata_reg_20,
	wrdata_reg_21,
	wrdata_reg_22,
	wrdata_reg_23,
	wrdata_reg_24,
	wrdata_reg_25,
	wrdata_reg_26,
	wrdata_reg_27,
	wrdata_reg_28,
	wrdata_reg_29,
	wrdata_reg_30,
	wrdata_reg_31,
	wrdata_reg_32,
	wrdata_reg_33,
	wrdata_reg_34,
	wrdata_reg_35,
	wrdata_reg_36,
	wrdata_reg_37,
	wrdata_reg_38,
	wrdata_reg_39,
	wrdata_reg_40,
	wrdata_reg_41,
	wrdata_reg_42,
	wrdata_reg_43,
	wrdata_reg_44,
	wrdata_reg_45,
	wrdata_reg_46,
	wrdata_reg_47,
	wrreq_reg1,
	avalon_streaming_sink_data,
	reset_sink_reset,
	avalon_streaming_sink_valid,
	clock_sink_clk)/* synthesis synthesis_greybox=0 */;
output 	wrdata_reg_0;
output 	wrdata_reg_1;
output 	wrdata_reg_2;
output 	wrdata_reg_3;
output 	wrdata_reg_4;
output 	wrdata_reg_5;
output 	wrdata_reg_6;
output 	wrdata_reg_7;
output 	wrdata_reg_8;
output 	wrdata_reg_9;
output 	wrdata_reg_10;
output 	wrdata_reg_11;
output 	wrdata_reg_12;
output 	wrdata_reg_13;
output 	wrdata_reg_14;
output 	wrdata_reg_15;
output 	wrdata_reg_16;
output 	wrdata_reg_17;
output 	wrdata_reg_18;
output 	wrdata_reg_19;
output 	wrdata_reg_20;
output 	wrdata_reg_21;
output 	wrdata_reg_22;
output 	wrdata_reg_23;
output 	wrdata_reg_24;
output 	wrdata_reg_25;
output 	wrdata_reg_26;
output 	wrdata_reg_27;
output 	wrdata_reg_28;
output 	wrdata_reg_29;
output 	wrdata_reg_30;
output 	wrdata_reg_31;
output 	wrdata_reg_32;
output 	wrdata_reg_33;
output 	wrdata_reg_34;
output 	wrdata_reg_35;
output 	wrdata_reg_36;
output 	wrdata_reg_37;
output 	wrdata_reg_38;
output 	wrdata_reg_39;
output 	wrdata_reg_40;
output 	wrdata_reg_41;
output 	wrdata_reg_42;
output 	wrdata_reg_43;
output 	wrdata_reg_44;
output 	wrdata_reg_45;
output 	wrdata_reg_46;
output 	wrdata_reg_47;
output 	wrreq_reg1;
input 	[47:0] avalon_streaming_sink_data;
input 	reset_sink_reset;
input 	avalon_streaming_sink_valid;
input 	clock_sink_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \wrdata_reg[0] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[0]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_0),
	.prn(vcc));
defparam \wrdata_reg[0] .is_wysiwyg = "true";
defparam \wrdata_reg[0] .power_up = "low";

dffeas \wrdata_reg[1] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[1]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_1),
	.prn(vcc));
defparam \wrdata_reg[1] .is_wysiwyg = "true";
defparam \wrdata_reg[1] .power_up = "low";

dffeas \wrdata_reg[2] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[2]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_2),
	.prn(vcc));
defparam \wrdata_reg[2] .is_wysiwyg = "true";
defparam \wrdata_reg[2] .power_up = "low";

dffeas \wrdata_reg[3] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[3]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_3),
	.prn(vcc));
defparam \wrdata_reg[3] .is_wysiwyg = "true";
defparam \wrdata_reg[3] .power_up = "low";

dffeas \wrdata_reg[4] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[4]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_4),
	.prn(vcc));
defparam \wrdata_reg[4] .is_wysiwyg = "true";
defparam \wrdata_reg[4] .power_up = "low";

dffeas \wrdata_reg[5] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[5]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_5),
	.prn(vcc));
defparam \wrdata_reg[5] .is_wysiwyg = "true";
defparam \wrdata_reg[5] .power_up = "low";

dffeas \wrdata_reg[6] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[6]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_6),
	.prn(vcc));
defparam \wrdata_reg[6] .is_wysiwyg = "true";
defparam \wrdata_reg[6] .power_up = "low";

dffeas \wrdata_reg[7] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[7]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_7),
	.prn(vcc));
defparam \wrdata_reg[7] .is_wysiwyg = "true";
defparam \wrdata_reg[7] .power_up = "low";

dffeas \wrdata_reg[8] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[8]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_8),
	.prn(vcc));
defparam \wrdata_reg[8] .is_wysiwyg = "true";
defparam \wrdata_reg[8] .power_up = "low";

dffeas \wrdata_reg[9] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[9]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_9),
	.prn(vcc));
defparam \wrdata_reg[9] .is_wysiwyg = "true";
defparam \wrdata_reg[9] .power_up = "low";

dffeas \wrdata_reg[10] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[10]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_10),
	.prn(vcc));
defparam \wrdata_reg[10] .is_wysiwyg = "true";
defparam \wrdata_reg[10] .power_up = "low";

dffeas \wrdata_reg[11] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[11]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_11),
	.prn(vcc));
defparam \wrdata_reg[11] .is_wysiwyg = "true";
defparam \wrdata_reg[11] .power_up = "low";

dffeas \wrdata_reg[12] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[12]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_12),
	.prn(vcc));
defparam \wrdata_reg[12] .is_wysiwyg = "true";
defparam \wrdata_reg[12] .power_up = "low";

dffeas \wrdata_reg[13] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[13]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_13),
	.prn(vcc));
defparam \wrdata_reg[13] .is_wysiwyg = "true";
defparam \wrdata_reg[13] .power_up = "low";

dffeas \wrdata_reg[14] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[14]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_14),
	.prn(vcc));
defparam \wrdata_reg[14] .is_wysiwyg = "true";
defparam \wrdata_reg[14] .power_up = "low";

dffeas \wrdata_reg[15] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[15]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_15),
	.prn(vcc));
defparam \wrdata_reg[15] .is_wysiwyg = "true";
defparam \wrdata_reg[15] .power_up = "low";

dffeas \wrdata_reg[16] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[16]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_16),
	.prn(vcc));
defparam \wrdata_reg[16] .is_wysiwyg = "true";
defparam \wrdata_reg[16] .power_up = "low";

dffeas \wrdata_reg[17] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[17]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_17),
	.prn(vcc));
defparam \wrdata_reg[17] .is_wysiwyg = "true";
defparam \wrdata_reg[17] .power_up = "low";

dffeas \wrdata_reg[18] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[18]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_18),
	.prn(vcc));
defparam \wrdata_reg[18] .is_wysiwyg = "true";
defparam \wrdata_reg[18] .power_up = "low";

dffeas \wrdata_reg[19] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[19]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_19),
	.prn(vcc));
defparam \wrdata_reg[19] .is_wysiwyg = "true";
defparam \wrdata_reg[19] .power_up = "low";

dffeas \wrdata_reg[20] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[20]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_20),
	.prn(vcc));
defparam \wrdata_reg[20] .is_wysiwyg = "true";
defparam \wrdata_reg[20] .power_up = "low";

dffeas \wrdata_reg[21] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[21]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_21),
	.prn(vcc));
defparam \wrdata_reg[21] .is_wysiwyg = "true";
defparam \wrdata_reg[21] .power_up = "low";

dffeas \wrdata_reg[22] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[22]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_22),
	.prn(vcc));
defparam \wrdata_reg[22] .is_wysiwyg = "true";
defparam \wrdata_reg[22] .power_up = "low";

dffeas \wrdata_reg[23] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[23]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_23),
	.prn(vcc));
defparam \wrdata_reg[23] .is_wysiwyg = "true";
defparam \wrdata_reg[23] .power_up = "low";

dffeas \wrdata_reg[24] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[24]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_24),
	.prn(vcc));
defparam \wrdata_reg[24] .is_wysiwyg = "true";
defparam \wrdata_reg[24] .power_up = "low";

dffeas \wrdata_reg[25] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[25]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_25),
	.prn(vcc));
defparam \wrdata_reg[25] .is_wysiwyg = "true";
defparam \wrdata_reg[25] .power_up = "low";

dffeas \wrdata_reg[26] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[26]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_26),
	.prn(vcc));
defparam \wrdata_reg[26] .is_wysiwyg = "true";
defparam \wrdata_reg[26] .power_up = "low";

dffeas \wrdata_reg[27] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[27]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_27),
	.prn(vcc));
defparam \wrdata_reg[27] .is_wysiwyg = "true";
defparam \wrdata_reg[27] .power_up = "low";

dffeas \wrdata_reg[28] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[28]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_28),
	.prn(vcc));
defparam \wrdata_reg[28] .is_wysiwyg = "true";
defparam \wrdata_reg[28] .power_up = "low";

dffeas \wrdata_reg[29] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[29]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_29),
	.prn(vcc));
defparam \wrdata_reg[29] .is_wysiwyg = "true";
defparam \wrdata_reg[29] .power_up = "low";

dffeas \wrdata_reg[30] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[30]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_30),
	.prn(vcc));
defparam \wrdata_reg[30] .is_wysiwyg = "true";
defparam \wrdata_reg[30] .power_up = "low";

dffeas \wrdata_reg[31] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[31]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_31),
	.prn(vcc));
defparam \wrdata_reg[31] .is_wysiwyg = "true";
defparam \wrdata_reg[31] .power_up = "low";

dffeas \wrdata_reg[32] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[32]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_32),
	.prn(vcc));
defparam \wrdata_reg[32] .is_wysiwyg = "true";
defparam \wrdata_reg[32] .power_up = "low";

dffeas \wrdata_reg[33] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[33]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_33),
	.prn(vcc));
defparam \wrdata_reg[33] .is_wysiwyg = "true";
defparam \wrdata_reg[33] .power_up = "low";

dffeas \wrdata_reg[34] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[34]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_34),
	.prn(vcc));
defparam \wrdata_reg[34] .is_wysiwyg = "true";
defparam \wrdata_reg[34] .power_up = "low";

dffeas \wrdata_reg[35] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[35]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_35),
	.prn(vcc));
defparam \wrdata_reg[35] .is_wysiwyg = "true";
defparam \wrdata_reg[35] .power_up = "low";

dffeas \wrdata_reg[36] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[36]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_36),
	.prn(vcc));
defparam \wrdata_reg[36] .is_wysiwyg = "true";
defparam \wrdata_reg[36] .power_up = "low";

dffeas \wrdata_reg[37] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[37]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_37),
	.prn(vcc));
defparam \wrdata_reg[37] .is_wysiwyg = "true";
defparam \wrdata_reg[37] .power_up = "low";

dffeas \wrdata_reg[38] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[38]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_38),
	.prn(vcc));
defparam \wrdata_reg[38] .is_wysiwyg = "true";
defparam \wrdata_reg[38] .power_up = "low";

dffeas \wrdata_reg[39] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[39]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_39),
	.prn(vcc));
defparam \wrdata_reg[39] .is_wysiwyg = "true";
defparam \wrdata_reg[39] .power_up = "low";

dffeas \wrdata_reg[40] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[40]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_40),
	.prn(vcc));
defparam \wrdata_reg[40] .is_wysiwyg = "true";
defparam \wrdata_reg[40] .power_up = "low";

dffeas \wrdata_reg[41] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[41]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_41),
	.prn(vcc));
defparam \wrdata_reg[41] .is_wysiwyg = "true";
defparam \wrdata_reg[41] .power_up = "low";

dffeas \wrdata_reg[42] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[42]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_42),
	.prn(vcc));
defparam \wrdata_reg[42] .is_wysiwyg = "true";
defparam \wrdata_reg[42] .power_up = "low";

dffeas \wrdata_reg[43] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[43]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_43),
	.prn(vcc));
defparam \wrdata_reg[43] .is_wysiwyg = "true";
defparam \wrdata_reg[43] .power_up = "low";

dffeas \wrdata_reg[44] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[44]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_44),
	.prn(vcc));
defparam \wrdata_reg[44] .is_wysiwyg = "true";
defparam \wrdata_reg[44] .power_up = "low";

dffeas \wrdata_reg[45] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[45]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_45),
	.prn(vcc));
defparam \wrdata_reg[45] .is_wysiwyg = "true";
defparam \wrdata_reg[45] .power_up = "low";

dffeas \wrdata_reg[46] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[46]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_46),
	.prn(vcc));
defparam \wrdata_reg[46] .is_wysiwyg = "true";
defparam \wrdata_reg[46] .power_up = "low";

dffeas \wrdata_reg[47] (
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_data[47]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrdata_reg_47),
	.prn(vcc));
defparam \wrdata_reg[47] .is_wysiwyg = "true";
defparam \wrdata_reg[47] .power_up = "low";

dffeas wrreq_reg(
	.clk(clock_sink_clk),
	.d(avalon_streaming_sink_valid),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wrreq_reg1),
	.prn(vcc));
defparam wrreq_reg.is_wysiwyg = "true";
defparam wrreq_reg.power_up = "low";

endmodule

module lms_dsp_fifo2avs (
	reset_sink_reset,
	valid_reg1,
	data_reg_21,
	data_reg_45,
	data_reg_20,
	data_reg_44,
	data_reg_19,
	data_reg_43,
	data_reg_18,
	data_reg_42,
	data_reg_17,
	data_reg_41,
	data_reg_16,
	data_reg_40,
	data_reg_15,
	data_reg_39,
	data_reg_14,
	data_reg_38,
	data_reg_12,
	data_reg_36,
	data_reg_13,
	data_reg_37,
	data_reg_9,
	data_reg_33,
	data_reg_8,
	data_reg_32,
	data_reg_7,
	data_reg_31,
	data_reg_6,
	data_reg_30,
	data_reg_5,
	data_reg_29,
	data_reg_4,
	data_reg_28,
	data_reg_3,
	data_reg_27,
	data_reg_2,
	data_reg_26,
	data_reg_0,
	data_reg_24,
	data_reg_1,
	data_reg_25,
	data_reg_11,
	data_reg_35,
	data_reg_10,
	data_reg_34,
	data_reg_23,
	data_reg_47,
	data_reg_22,
	data_reg_46,
	clock_sink_clk,
	fifo_wrreq,
	fifo_wdata)/* synthesis synthesis_greybox=0 */;
input 	reset_sink_reset;
output 	valid_reg1;
output 	data_reg_21;
output 	data_reg_45;
output 	data_reg_20;
output 	data_reg_44;
output 	data_reg_19;
output 	data_reg_43;
output 	data_reg_18;
output 	data_reg_42;
output 	data_reg_17;
output 	data_reg_41;
output 	data_reg_16;
output 	data_reg_40;
output 	data_reg_15;
output 	data_reg_39;
output 	data_reg_14;
output 	data_reg_38;
output 	data_reg_12;
output 	data_reg_36;
output 	data_reg_13;
output 	data_reg_37;
output 	data_reg_9;
output 	data_reg_33;
output 	data_reg_8;
output 	data_reg_32;
output 	data_reg_7;
output 	data_reg_31;
output 	data_reg_6;
output 	data_reg_30;
output 	data_reg_5;
output 	data_reg_29;
output 	data_reg_4;
output 	data_reg_28;
output 	data_reg_3;
output 	data_reg_27;
output 	data_reg_2;
output 	data_reg_26;
output 	data_reg_0;
output 	data_reg_24;
output 	data_reg_1;
output 	data_reg_25;
output 	data_reg_11;
output 	data_reg_35;
output 	data_reg_10;
output 	data_reg_34;
output 	data_reg_23;
output 	data_reg_47;
output 	data_reg_22;
output 	data_reg_46;
input 	clock_sink_clk;
input 	fifo_wrreq;
input 	[47:0] fifo_wdata;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas valid_reg(
	.clk(clock_sink_clk),
	.d(fifo_wrreq),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(valid_reg1),
	.prn(vcc));
defparam valid_reg.is_wysiwyg = "true";
defparam valid_reg.power_up = "low";

dffeas \data_reg[21] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[21]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_21),
	.prn(vcc));
defparam \data_reg[21] .is_wysiwyg = "true";
defparam \data_reg[21] .power_up = "low";

dffeas \data_reg[45] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[45]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_45),
	.prn(vcc));
defparam \data_reg[45] .is_wysiwyg = "true";
defparam \data_reg[45] .power_up = "low";

dffeas \data_reg[20] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[20]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_20),
	.prn(vcc));
defparam \data_reg[20] .is_wysiwyg = "true";
defparam \data_reg[20] .power_up = "low";

dffeas \data_reg[44] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[44]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_44),
	.prn(vcc));
defparam \data_reg[44] .is_wysiwyg = "true";
defparam \data_reg[44] .power_up = "low";

dffeas \data_reg[19] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[19]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_19),
	.prn(vcc));
defparam \data_reg[19] .is_wysiwyg = "true";
defparam \data_reg[19] .power_up = "low";

dffeas \data_reg[43] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[43]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_43),
	.prn(vcc));
defparam \data_reg[43] .is_wysiwyg = "true";
defparam \data_reg[43] .power_up = "low";

dffeas \data_reg[18] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[18]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_18),
	.prn(vcc));
defparam \data_reg[18] .is_wysiwyg = "true";
defparam \data_reg[18] .power_up = "low";

dffeas \data_reg[42] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[42]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_42),
	.prn(vcc));
defparam \data_reg[42] .is_wysiwyg = "true";
defparam \data_reg[42] .power_up = "low";

dffeas \data_reg[17] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[17]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_17),
	.prn(vcc));
defparam \data_reg[17] .is_wysiwyg = "true";
defparam \data_reg[17] .power_up = "low";

dffeas \data_reg[41] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[41]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_41),
	.prn(vcc));
defparam \data_reg[41] .is_wysiwyg = "true";
defparam \data_reg[41] .power_up = "low";

dffeas \data_reg[16] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[16]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_16),
	.prn(vcc));
defparam \data_reg[16] .is_wysiwyg = "true";
defparam \data_reg[16] .power_up = "low";

dffeas \data_reg[40] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[40]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_40),
	.prn(vcc));
defparam \data_reg[40] .is_wysiwyg = "true";
defparam \data_reg[40] .power_up = "low";

dffeas \data_reg[15] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[15]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_15),
	.prn(vcc));
defparam \data_reg[15] .is_wysiwyg = "true";
defparam \data_reg[15] .power_up = "low";

dffeas \data_reg[39] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[39]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_39),
	.prn(vcc));
defparam \data_reg[39] .is_wysiwyg = "true";
defparam \data_reg[39] .power_up = "low";

dffeas \data_reg[14] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[14]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_14),
	.prn(vcc));
defparam \data_reg[14] .is_wysiwyg = "true";
defparam \data_reg[14] .power_up = "low";

dffeas \data_reg[38] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[38]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_38),
	.prn(vcc));
defparam \data_reg[38] .is_wysiwyg = "true";
defparam \data_reg[38] .power_up = "low";

dffeas \data_reg[12] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[12]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_12),
	.prn(vcc));
defparam \data_reg[12] .is_wysiwyg = "true";
defparam \data_reg[12] .power_up = "low";

dffeas \data_reg[36] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[36]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_36),
	.prn(vcc));
defparam \data_reg[36] .is_wysiwyg = "true";
defparam \data_reg[36] .power_up = "low";

dffeas \data_reg[13] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[13]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_13),
	.prn(vcc));
defparam \data_reg[13] .is_wysiwyg = "true";
defparam \data_reg[13] .power_up = "low";

dffeas \data_reg[37] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[37]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_37),
	.prn(vcc));
defparam \data_reg[37] .is_wysiwyg = "true";
defparam \data_reg[37] .power_up = "low";

dffeas \data_reg[9] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[9]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_9),
	.prn(vcc));
defparam \data_reg[9] .is_wysiwyg = "true";
defparam \data_reg[9] .power_up = "low";

dffeas \data_reg[33] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[33]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_33),
	.prn(vcc));
defparam \data_reg[33] .is_wysiwyg = "true";
defparam \data_reg[33] .power_up = "low";

dffeas \data_reg[8] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[8]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_8),
	.prn(vcc));
defparam \data_reg[8] .is_wysiwyg = "true";
defparam \data_reg[8] .power_up = "low";

dffeas \data_reg[32] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[32]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_32),
	.prn(vcc));
defparam \data_reg[32] .is_wysiwyg = "true";
defparam \data_reg[32] .power_up = "low";

dffeas \data_reg[7] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[7]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_7),
	.prn(vcc));
defparam \data_reg[7] .is_wysiwyg = "true";
defparam \data_reg[7] .power_up = "low";

dffeas \data_reg[31] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[31]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_31),
	.prn(vcc));
defparam \data_reg[31] .is_wysiwyg = "true";
defparam \data_reg[31] .power_up = "low";

dffeas \data_reg[6] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[6]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_6),
	.prn(vcc));
defparam \data_reg[6] .is_wysiwyg = "true";
defparam \data_reg[6] .power_up = "low";

dffeas \data_reg[30] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[30]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_30),
	.prn(vcc));
defparam \data_reg[30] .is_wysiwyg = "true";
defparam \data_reg[30] .power_up = "low";

dffeas \data_reg[5] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[5]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_5),
	.prn(vcc));
defparam \data_reg[5] .is_wysiwyg = "true";
defparam \data_reg[5] .power_up = "low";

dffeas \data_reg[29] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[29]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_29),
	.prn(vcc));
defparam \data_reg[29] .is_wysiwyg = "true";
defparam \data_reg[29] .power_up = "low";

dffeas \data_reg[4] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[4]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_4),
	.prn(vcc));
defparam \data_reg[4] .is_wysiwyg = "true";
defparam \data_reg[4] .power_up = "low";

dffeas \data_reg[28] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[28]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_28),
	.prn(vcc));
defparam \data_reg[28] .is_wysiwyg = "true";
defparam \data_reg[28] .power_up = "low";

dffeas \data_reg[3] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[3]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_3),
	.prn(vcc));
defparam \data_reg[3] .is_wysiwyg = "true";
defparam \data_reg[3] .power_up = "low";

dffeas \data_reg[27] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[27]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_27),
	.prn(vcc));
defparam \data_reg[27] .is_wysiwyg = "true";
defparam \data_reg[27] .power_up = "low";

dffeas \data_reg[2] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[2]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_2),
	.prn(vcc));
defparam \data_reg[2] .is_wysiwyg = "true";
defparam \data_reg[2] .power_up = "low";

dffeas \data_reg[26] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[26]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_26),
	.prn(vcc));
defparam \data_reg[26] .is_wysiwyg = "true";
defparam \data_reg[26] .power_up = "low";

dffeas \data_reg[0] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[0]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_0),
	.prn(vcc));
defparam \data_reg[0] .is_wysiwyg = "true";
defparam \data_reg[0] .power_up = "low";

dffeas \data_reg[24] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[24]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_24),
	.prn(vcc));
defparam \data_reg[24] .is_wysiwyg = "true";
defparam \data_reg[24] .power_up = "low";

dffeas \data_reg[1] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[1]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_1),
	.prn(vcc));
defparam \data_reg[1] .is_wysiwyg = "true";
defparam \data_reg[1] .power_up = "low";

dffeas \data_reg[25] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[25]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_25),
	.prn(vcc));
defparam \data_reg[25] .is_wysiwyg = "true";
defparam \data_reg[25] .power_up = "low";

dffeas \data_reg[11] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[11]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_11),
	.prn(vcc));
defparam \data_reg[11] .is_wysiwyg = "true";
defparam \data_reg[11] .power_up = "low";

dffeas \data_reg[35] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[35]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_35),
	.prn(vcc));
defparam \data_reg[35] .is_wysiwyg = "true";
defparam \data_reg[35] .power_up = "low";

dffeas \data_reg[10] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[10]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_10),
	.prn(vcc));
defparam \data_reg[10] .is_wysiwyg = "true";
defparam \data_reg[10] .power_up = "low";

dffeas \data_reg[34] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[34]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_34),
	.prn(vcc));
defparam \data_reg[34] .is_wysiwyg = "true";
defparam \data_reg[34] .power_up = "low";

dffeas \data_reg[23] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[23]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_23),
	.prn(vcc));
defparam \data_reg[23] .is_wysiwyg = "true";
defparam \data_reg[23] .power_up = "low";

dffeas \data_reg[47] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[47]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_47),
	.prn(vcc));
defparam \data_reg[47] .is_wysiwyg = "true";
defparam \data_reg[47] .power_up = "low";

dffeas \data_reg[22] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[22]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_22),
	.prn(vcc));
defparam \data_reg[22] .is_wysiwyg = "true";
defparam \data_reg[22] .power_up = "low";

dffeas \data_reg[46] (
	.clk(clock_sink_clk),
	.d(fifo_wdata[46]),
	.asdata(vcc),
	.clrn(reset_sink_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_reg_46),
	.prn(vcc));
defparam \data_reg[46] .is_wysiwyg = "true";
defparam \data_reg[46] .power_up = "low";

endmodule

module lms_dsp_lms_dsp_avalon_st_adapter (
	out_data_0,
	altera_reset_synchronizer_int_chain_out,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_5,
	out_data_6,
	out_data_7,
	out_data_8,
	out_data_9,
	out_data_10,
	out_data_11,
	out_data_12,
	out_data_13,
	out_data_14,
	out_data_15,
	out_data_16,
	out_data_17,
	out_data_18,
	out_data_19,
	out_data_20,
	out_data_21,
	out_data_22,
	out_data_23,
	out_data_24,
	out_data_25,
	out_data_26,
	out_data_27,
	out_data_28,
	out_data_29,
	out_data_30,
	out_data_31,
	out_data_32,
	out_data_33,
	out_data_34,
	out_data_35,
	out_data_36,
	out_data_37,
	out_data_38,
	out_data_39,
	out_data_40,
	out_data_41,
	out_data_42,
	out_data_43,
	out_data_44,
	out_data_45,
	out_data_46,
	out_data_47,
	out_valid,
	avalon_streaming_source_data_0,
	avalon_streaming_source_data_1,
	avalon_streaming_source_data_2,
	avalon_streaming_source_data_3,
	avalon_streaming_source_data_4,
	avalon_streaming_source_data_5,
	avalon_streaming_source_data_6,
	avalon_streaming_source_data_7,
	avalon_streaming_source_data_8,
	avalon_streaming_source_data_9,
	avalon_streaming_source_data_10,
	avalon_streaming_source_data_11,
	avalon_streaming_source_data_12,
	avalon_streaming_source_data_13,
	avalon_streaming_source_data_14,
	avalon_streaming_source_data_15,
	avalon_streaming_source_data_16,
	avalon_streaming_source_data_17,
	avalon_streaming_source_data_18,
	avalon_streaming_source_data_19,
	avalon_streaming_source_data_20,
	avalon_streaming_source_data_21,
	avalon_streaming_source_data_22,
	avalon_streaming_source_data_23,
	delay_reg_24_3,
	clk_clk)/* synthesis synthesis_greybox=0 */;
output 	out_data_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	out_data_1;
output 	out_data_2;
output 	out_data_3;
output 	out_data_4;
output 	out_data_5;
output 	out_data_6;
output 	out_data_7;
output 	out_data_8;
output 	out_data_9;
output 	out_data_10;
output 	out_data_11;
output 	out_data_12;
output 	out_data_13;
output 	out_data_14;
output 	out_data_15;
output 	out_data_16;
output 	out_data_17;
output 	out_data_18;
output 	out_data_19;
output 	out_data_20;
output 	out_data_21;
output 	out_data_22;
output 	out_data_23;
output 	out_data_24;
output 	out_data_25;
output 	out_data_26;
output 	out_data_27;
output 	out_data_28;
output 	out_data_29;
output 	out_data_30;
output 	out_data_31;
output 	out_data_32;
output 	out_data_33;
output 	out_data_34;
output 	out_data_35;
output 	out_data_36;
output 	out_data_37;
output 	out_data_38;
output 	out_data_39;
output 	out_data_40;
output 	out_data_41;
output 	out_data_42;
output 	out_data_43;
output 	out_data_44;
output 	out_data_45;
output 	out_data_46;
output 	out_data_47;
output 	out_valid;
input 	avalon_streaming_source_data_0;
input 	avalon_streaming_source_data_1;
input 	avalon_streaming_source_data_2;
input 	avalon_streaming_source_data_3;
input 	avalon_streaming_source_data_4;
input 	avalon_streaming_source_data_5;
input 	avalon_streaming_source_data_6;
input 	avalon_streaming_source_data_7;
input 	avalon_streaming_source_data_8;
input 	avalon_streaming_source_data_9;
input 	avalon_streaming_source_data_10;
input 	avalon_streaming_source_data_11;
input 	avalon_streaming_source_data_12;
input 	avalon_streaming_source_data_13;
input 	avalon_streaming_source_data_14;
input 	avalon_streaming_source_data_15;
input 	avalon_streaming_source_data_16;
input 	avalon_streaming_source_data_17;
input 	avalon_streaming_source_data_18;
input 	avalon_streaming_source_data_19;
input 	avalon_streaming_source_data_20;
input 	avalon_streaming_source_data_21;
input 	avalon_streaming_source_data_22;
input 	avalon_streaming_source_data_23;
input 	delay_reg_24_3;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



lms_dsp_lms_dsp_avalon_st_adapter_data_format_adapter_0 data_format_adapter_0(
	.out_data_0(out_data_0),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.out_data_1(out_data_1),
	.out_data_2(out_data_2),
	.out_data_3(out_data_3),
	.out_data_4(out_data_4),
	.out_data_5(out_data_5),
	.out_data_6(out_data_6),
	.out_data_7(out_data_7),
	.out_data_8(out_data_8),
	.out_data_9(out_data_9),
	.out_data_10(out_data_10),
	.out_data_11(out_data_11),
	.out_data_12(out_data_12),
	.out_data_13(out_data_13),
	.out_data_14(out_data_14),
	.out_data_15(out_data_15),
	.out_data_16(out_data_16),
	.out_data_17(out_data_17),
	.out_data_18(out_data_18),
	.out_data_19(out_data_19),
	.out_data_20(out_data_20),
	.out_data_21(out_data_21),
	.out_data_22(out_data_22),
	.out_data_23(out_data_23),
	.out_data_24(out_data_24),
	.out_data_25(out_data_25),
	.out_data_26(out_data_26),
	.out_data_27(out_data_27),
	.out_data_28(out_data_28),
	.out_data_29(out_data_29),
	.out_data_30(out_data_30),
	.out_data_31(out_data_31),
	.out_data_32(out_data_32),
	.out_data_33(out_data_33),
	.out_data_34(out_data_34),
	.out_data_35(out_data_35),
	.out_data_36(out_data_36),
	.out_data_37(out_data_37),
	.out_data_38(out_data_38),
	.out_data_39(out_data_39),
	.out_data_40(out_data_40),
	.out_data_41(out_data_41),
	.out_data_42(out_data_42),
	.out_data_43(out_data_43),
	.out_data_44(out_data_44),
	.out_data_45(out_data_45),
	.out_data_46(out_data_46),
	.out_data_47(out_data_47),
	.out_valid1(out_valid),
	.in_data({avalon_streaming_source_data_23,avalon_streaming_source_data_22,avalon_streaming_source_data_21,avalon_streaming_source_data_20,avalon_streaming_source_data_19,avalon_streaming_source_data_18,avalon_streaming_source_data_17,avalon_streaming_source_data_16,
avalon_streaming_source_data_15,avalon_streaming_source_data_14,avalon_streaming_source_data_13,avalon_streaming_source_data_12,avalon_streaming_source_data_11,avalon_streaming_source_data_10,avalon_streaming_source_data_9,avalon_streaming_source_data_8,
avalon_streaming_source_data_7,avalon_streaming_source_data_6,avalon_streaming_source_data_5,avalon_streaming_source_data_4,avalon_streaming_source_data_3,avalon_streaming_source_data_2,avalon_streaming_source_data_1,avalon_streaming_source_data_0}),
	.in_valid(delay_reg_24_3),
	.clk(clk_clk));

endmodule

module lms_dsp_lms_dsp_avalon_st_adapter_data_format_adapter_0 (
	out_data_0,
	reset_n,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_5,
	out_data_6,
	out_data_7,
	out_data_8,
	out_data_9,
	out_data_10,
	out_data_11,
	out_data_12,
	out_data_13,
	out_data_14,
	out_data_15,
	out_data_16,
	out_data_17,
	out_data_18,
	out_data_19,
	out_data_20,
	out_data_21,
	out_data_22,
	out_data_23,
	out_data_24,
	out_data_25,
	out_data_26,
	out_data_27,
	out_data_28,
	out_data_29,
	out_data_30,
	out_data_31,
	out_data_32,
	out_data_33,
	out_data_34,
	out_data_35,
	out_data_36,
	out_data_37,
	out_data_38,
	out_data_39,
	out_data_40,
	out_data_41,
	out_data_42,
	out_data_43,
	out_data_44,
	out_data_45,
	out_data_46,
	out_data_47,
	out_valid1,
	in_data,
	in_valid,
	clk)/* synthesis synthesis_greybox=0 */;
output 	out_data_0;
input 	reset_n;
output 	out_data_1;
output 	out_data_2;
output 	out_data_3;
output 	out_data_4;
output 	out_data_5;
output 	out_data_6;
output 	out_data_7;
output 	out_data_8;
output 	out_data_9;
output 	out_data_10;
output 	out_data_11;
output 	out_data_12;
output 	out_data_13;
output 	out_data_14;
output 	out_data_15;
output 	out_data_16;
output 	out_data_17;
output 	out_data_18;
output 	out_data_19;
output 	out_data_20;
output 	out_data_21;
output 	out_data_22;
output 	out_data_23;
output 	out_data_24;
output 	out_data_25;
output 	out_data_26;
output 	out_data_27;
output 	out_data_28;
output 	out_data_29;
output 	out_data_30;
output 	out_data_31;
output 	out_data_32;
output 	out_data_33;
output 	out_data_34;
output 	out_data_35;
output 	out_data_36;
output 	out_data_37;
output 	out_data_38;
output 	out_data_39;
output 	out_data_40;
output 	out_data_41;
output 	out_data_42;
output 	out_data_43;
output 	out_data_44;
output 	out_data_45;
output 	out_data_46;
output 	out_data_47;
output 	out_valid1;
input 	[23:0] in_data;
input 	in_valid;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a_data1[0]~q ;
wire \in_ready_d1~q ;
wire \state[0]~0_combout ;
wire \state_d1[0]~q ;
wire \a_valid~q ;
wire \Mux2~0_combout ;
wire \state_register[0]~q ;
wire \b_data[0]~0_combout ;
wire \a_data1[1]~q ;
wire \b_data[1]~1_combout ;
wire \a_data1[2]~q ;
wire \b_data[2]~2_combout ;
wire \a_data1[3]~q ;
wire \b_data[3]~3_combout ;
wire \a_data1[4]~q ;
wire \b_data[4]~4_combout ;
wire \a_data1[5]~q ;
wire \b_data[5]~5_combout ;
wire \a_data1[6]~q ;
wire \b_data[6]~6_combout ;
wire \a_data1[7]~q ;
wire \b_data[7]~7_combout ;
wire \a_data1[8]~q ;
wire \b_data[8]~8_combout ;
wire \a_data1[9]~q ;
wire \b_data[9]~9_combout ;
wire \a_data1[10]~q ;
wire \b_data[10]~10_combout ;
wire \a_data1[11]~q ;
wire \b_data[11]~11_combout ;
wire \a_data0[0]~q ;
wire \b_data[12]~12_combout ;
wire \a_data0[1]~q ;
wire \b_data[13]~13_combout ;
wire \a_data0[2]~q ;
wire \b_data[14]~14_combout ;
wire \a_data0[3]~q ;
wire \b_data[15]~15_combout ;
wire \a_data0[4]~q ;
wire \b_data[16]~16_combout ;
wire \a_data0[5]~q ;
wire \b_data[17]~17_combout ;
wire \a_data0[6]~q ;
wire \b_data[18]~18_combout ;
wire \a_data0[7]~q ;
wire \b_data[19]~19_combout ;
wire \a_data0[8]~q ;
wire \b_data[20]~20_combout ;
wire \a_data0[9]~q ;
wire \b_data[21]~21_combout ;
wire \a_data0[10]~q ;
wire \b_data[22]~22_combout ;
wire \a_data0[11]~q ;
wire \b_data[23]~23_combout ;
wire \Mux5~0_combout ;
wire \data1_register[0]~q ;
wire \b_data[24]~24_combout ;
wire \data1_register[1]~q ;
wire \b_data[25]~25_combout ;
wire \data1_register[2]~q ;
wire \b_data[26]~26_combout ;
wire \data1_register[3]~q ;
wire \b_data[27]~27_combout ;
wire \data1_register[4]~q ;
wire \b_data[28]~28_combout ;
wire \data1_register[5]~q ;
wire \b_data[29]~29_combout ;
wire \data1_register[6]~q ;
wire \b_data[30]~30_combout ;
wire \data1_register[7]~q ;
wire \b_data[31]~31_combout ;
wire \data1_register[8]~q ;
wire \b_data[32]~32_combout ;
wire \data1_register[9]~q ;
wire \b_data[33]~33_combout ;
wire \data1_register[10]~q ;
wire \b_data[34]~34_combout ;
wire \data1_register[11]~q ;
wire \b_data[35]~35_combout ;
wire \data0_register[0]~q ;
wire \b_data[36]~36_combout ;
wire \data0_register[1]~q ;
wire \b_data[37]~37_combout ;
wire \data0_register[2]~q ;
wire \b_data[38]~38_combout ;
wire \data0_register[3]~q ;
wire \b_data[39]~39_combout ;
wire \data0_register[4]~q ;
wire \b_data[40]~40_combout ;
wire \data0_register[5]~q ;
wire \b_data[41]~41_combout ;
wire \data0_register[6]~q ;
wire \b_data[42]~42_combout ;
wire \data0_register[7]~q ;
wire \b_data[43]~43_combout ;
wire \data0_register[8]~q ;
wire \b_data[44]~44_combout ;
wire \data0_register[9]~q ;
wire \b_data[45]~45_combout ;
wire \data0_register[10]~q ;
wire \b_data[46]~46_combout ;
wire \data0_register[11]~q ;
wire \b_data[47]~47_combout ;
wire \Mux3~0_combout ;


dffeas \out_data[0] (
	.clk(clk),
	.d(\b_data[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_0),
	.prn(vcc));
defparam \out_data[0] .is_wysiwyg = "true";
defparam \out_data[0] .power_up = "low";

dffeas \out_data[1] (
	.clk(clk),
	.d(\b_data[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_1),
	.prn(vcc));
defparam \out_data[1] .is_wysiwyg = "true";
defparam \out_data[1] .power_up = "low";

dffeas \out_data[2] (
	.clk(clk),
	.d(\b_data[2]~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_2),
	.prn(vcc));
defparam \out_data[2] .is_wysiwyg = "true";
defparam \out_data[2] .power_up = "low";

dffeas \out_data[3] (
	.clk(clk),
	.d(\b_data[3]~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_3),
	.prn(vcc));
defparam \out_data[3] .is_wysiwyg = "true";
defparam \out_data[3] .power_up = "low";

dffeas \out_data[4] (
	.clk(clk),
	.d(\b_data[4]~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_4),
	.prn(vcc));
defparam \out_data[4] .is_wysiwyg = "true";
defparam \out_data[4] .power_up = "low";

dffeas \out_data[5] (
	.clk(clk),
	.d(\b_data[5]~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_5),
	.prn(vcc));
defparam \out_data[5] .is_wysiwyg = "true";
defparam \out_data[5] .power_up = "low";

dffeas \out_data[6] (
	.clk(clk),
	.d(\b_data[6]~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_6),
	.prn(vcc));
defparam \out_data[6] .is_wysiwyg = "true";
defparam \out_data[6] .power_up = "low";

dffeas \out_data[7] (
	.clk(clk),
	.d(\b_data[7]~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_7),
	.prn(vcc));
defparam \out_data[7] .is_wysiwyg = "true";
defparam \out_data[7] .power_up = "low";

dffeas \out_data[8] (
	.clk(clk),
	.d(\b_data[8]~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_8),
	.prn(vcc));
defparam \out_data[8] .is_wysiwyg = "true";
defparam \out_data[8] .power_up = "low";

dffeas \out_data[9] (
	.clk(clk),
	.d(\b_data[9]~9_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_9),
	.prn(vcc));
defparam \out_data[9] .is_wysiwyg = "true";
defparam \out_data[9] .power_up = "low";

dffeas \out_data[10] (
	.clk(clk),
	.d(\b_data[10]~10_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_10),
	.prn(vcc));
defparam \out_data[10] .is_wysiwyg = "true";
defparam \out_data[10] .power_up = "low";

dffeas \out_data[11] (
	.clk(clk),
	.d(\b_data[11]~11_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_11),
	.prn(vcc));
defparam \out_data[11] .is_wysiwyg = "true";
defparam \out_data[11] .power_up = "low";

dffeas \out_data[12] (
	.clk(clk),
	.d(\b_data[12]~12_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_12),
	.prn(vcc));
defparam \out_data[12] .is_wysiwyg = "true";
defparam \out_data[12] .power_up = "low";

dffeas \out_data[13] (
	.clk(clk),
	.d(\b_data[13]~13_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_13),
	.prn(vcc));
defparam \out_data[13] .is_wysiwyg = "true";
defparam \out_data[13] .power_up = "low";

dffeas \out_data[14] (
	.clk(clk),
	.d(\b_data[14]~14_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_14),
	.prn(vcc));
defparam \out_data[14] .is_wysiwyg = "true";
defparam \out_data[14] .power_up = "low";

dffeas \out_data[15] (
	.clk(clk),
	.d(\b_data[15]~15_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_15),
	.prn(vcc));
defparam \out_data[15] .is_wysiwyg = "true";
defparam \out_data[15] .power_up = "low";

dffeas \out_data[16] (
	.clk(clk),
	.d(\b_data[16]~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_16),
	.prn(vcc));
defparam \out_data[16] .is_wysiwyg = "true";
defparam \out_data[16] .power_up = "low";

dffeas \out_data[17] (
	.clk(clk),
	.d(\b_data[17]~17_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_17),
	.prn(vcc));
defparam \out_data[17] .is_wysiwyg = "true";
defparam \out_data[17] .power_up = "low";

dffeas \out_data[18] (
	.clk(clk),
	.d(\b_data[18]~18_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_18),
	.prn(vcc));
defparam \out_data[18] .is_wysiwyg = "true";
defparam \out_data[18] .power_up = "low";

dffeas \out_data[19] (
	.clk(clk),
	.d(\b_data[19]~19_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_19),
	.prn(vcc));
defparam \out_data[19] .is_wysiwyg = "true";
defparam \out_data[19] .power_up = "low";

dffeas \out_data[20] (
	.clk(clk),
	.d(\b_data[20]~20_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_20),
	.prn(vcc));
defparam \out_data[20] .is_wysiwyg = "true";
defparam \out_data[20] .power_up = "low";

dffeas \out_data[21] (
	.clk(clk),
	.d(\b_data[21]~21_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_21),
	.prn(vcc));
defparam \out_data[21] .is_wysiwyg = "true";
defparam \out_data[21] .power_up = "low";

dffeas \out_data[22] (
	.clk(clk),
	.d(\b_data[22]~22_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_22),
	.prn(vcc));
defparam \out_data[22] .is_wysiwyg = "true";
defparam \out_data[22] .power_up = "low";

dffeas \out_data[23] (
	.clk(clk),
	.d(\b_data[23]~23_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_23),
	.prn(vcc));
defparam \out_data[23] .is_wysiwyg = "true";
defparam \out_data[23] .power_up = "low";

dffeas \out_data[24] (
	.clk(clk),
	.d(\b_data[24]~24_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_24),
	.prn(vcc));
defparam \out_data[24] .is_wysiwyg = "true";
defparam \out_data[24] .power_up = "low";

dffeas \out_data[25] (
	.clk(clk),
	.d(\b_data[25]~25_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_25),
	.prn(vcc));
defparam \out_data[25] .is_wysiwyg = "true";
defparam \out_data[25] .power_up = "low";

dffeas \out_data[26] (
	.clk(clk),
	.d(\b_data[26]~26_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_26),
	.prn(vcc));
defparam \out_data[26] .is_wysiwyg = "true";
defparam \out_data[26] .power_up = "low";

dffeas \out_data[27] (
	.clk(clk),
	.d(\b_data[27]~27_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_27),
	.prn(vcc));
defparam \out_data[27] .is_wysiwyg = "true";
defparam \out_data[27] .power_up = "low";

dffeas \out_data[28] (
	.clk(clk),
	.d(\b_data[28]~28_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_28),
	.prn(vcc));
defparam \out_data[28] .is_wysiwyg = "true";
defparam \out_data[28] .power_up = "low";

dffeas \out_data[29] (
	.clk(clk),
	.d(\b_data[29]~29_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_29),
	.prn(vcc));
defparam \out_data[29] .is_wysiwyg = "true";
defparam \out_data[29] .power_up = "low";

dffeas \out_data[30] (
	.clk(clk),
	.d(\b_data[30]~30_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_30),
	.prn(vcc));
defparam \out_data[30] .is_wysiwyg = "true";
defparam \out_data[30] .power_up = "low";

dffeas \out_data[31] (
	.clk(clk),
	.d(\b_data[31]~31_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_31),
	.prn(vcc));
defparam \out_data[31] .is_wysiwyg = "true";
defparam \out_data[31] .power_up = "low";

dffeas \out_data[32] (
	.clk(clk),
	.d(\b_data[32]~32_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_32),
	.prn(vcc));
defparam \out_data[32] .is_wysiwyg = "true";
defparam \out_data[32] .power_up = "low";

dffeas \out_data[33] (
	.clk(clk),
	.d(\b_data[33]~33_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_33),
	.prn(vcc));
defparam \out_data[33] .is_wysiwyg = "true";
defparam \out_data[33] .power_up = "low";

dffeas \out_data[34] (
	.clk(clk),
	.d(\b_data[34]~34_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_34),
	.prn(vcc));
defparam \out_data[34] .is_wysiwyg = "true";
defparam \out_data[34] .power_up = "low";

dffeas \out_data[35] (
	.clk(clk),
	.d(\b_data[35]~35_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_35),
	.prn(vcc));
defparam \out_data[35] .is_wysiwyg = "true";
defparam \out_data[35] .power_up = "low";

dffeas \out_data[36] (
	.clk(clk),
	.d(\b_data[36]~36_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_36),
	.prn(vcc));
defparam \out_data[36] .is_wysiwyg = "true";
defparam \out_data[36] .power_up = "low";

dffeas \out_data[37] (
	.clk(clk),
	.d(\b_data[37]~37_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_37),
	.prn(vcc));
defparam \out_data[37] .is_wysiwyg = "true";
defparam \out_data[37] .power_up = "low";

dffeas \out_data[38] (
	.clk(clk),
	.d(\b_data[38]~38_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_38),
	.prn(vcc));
defparam \out_data[38] .is_wysiwyg = "true";
defparam \out_data[38] .power_up = "low";

dffeas \out_data[39] (
	.clk(clk),
	.d(\b_data[39]~39_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_39),
	.prn(vcc));
defparam \out_data[39] .is_wysiwyg = "true";
defparam \out_data[39] .power_up = "low";

dffeas \out_data[40] (
	.clk(clk),
	.d(\b_data[40]~40_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_40),
	.prn(vcc));
defparam \out_data[40] .is_wysiwyg = "true";
defparam \out_data[40] .power_up = "low";

dffeas \out_data[41] (
	.clk(clk),
	.d(\b_data[41]~41_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_41),
	.prn(vcc));
defparam \out_data[41] .is_wysiwyg = "true";
defparam \out_data[41] .power_up = "low";

dffeas \out_data[42] (
	.clk(clk),
	.d(\b_data[42]~42_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_42),
	.prn(vcc));
defparam \out_data[42] .is_wysiwyg = "true";
defparam \out_data[42] .power_up = "low";

dffeas \out_data[43] (
	.clk(clk),
	.d(\b_data[43]~43_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_43),
	.prn(vcc));
defparam \out_data[43] .is_wysiwyg = "true";
defparam \out_data[43] .power_up = "low";

dffeas \out_data[44] (
	.clk(clk),
	.d(\b_data[44]~44_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_44),
	.prn(vcc));
defparam \out_data[44] .is_wysiwyg = "true";
defparam \out_data[44] .power_up = "low";

dffeas \out_data[45] (
	.clk(clk),
	.d(\b_data[45]~45_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_45),
	.prn(vcc));
defparam \out_data[45] .is_wysiwyg = "true";
defparam \out_data[45] .power_up = "low";

dffeas \out_data[46] (
	.clk(clk),
	.d(\b_data[46]~46_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_46),
	.prn(vcc));
defparam \out_data[46] .is_wysiwyg = "true";
defparam \out_data[46] .power_up = "low";

dffeas \out_data[47] (
	.clk(clk),
	.d(\b_data[47]~47_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_47),
	.prn(vcc));
defparam \out_data[47] .is_wysiwyg = "true";
defparam \out_data[47] .power_up = "low";

dffeas out_valid(
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

dffeas \a_data1[0] (
	.clk(clk),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data1[0]~q ),
	.prn(vcc));
defparam \a_data1[0] .is_wysiwyg = "true";
defparam \a_data1[0] .power_up = "low";

dffeas in_ready_d1(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_ready_d1~q ),
	.prn(vcc));
defparam in_ready_d1.is_wysiwyg = "true";
defparam in_ready_d1.power_up = "low";

fiftyfivenm_lcell_comb \state[0]~0 (
	.dataa(\state_register[0]~q ),
	.datab(\state_d1[0]~q ),
	.datac(gnd),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\state[0]~0_combout ),
	.cout());
defparam \state[0]~0 .lut_mask = 16'hAACC;
defparam \state[0]~0 .sum_lutc_input = "datac";

dffeas \state_d1[0] (
	.clk(clk),
	.d(\state[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state_d1[0]~q ),
	.prn(vcc));
defparam \state_d1[0] .is_wysiwyg = "true";
defparam \state_d1[0] .power_up = "low";

dffeas a_valid(
	.clk(clk),
	.d(in_valid),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_valid~q ),
	.prn(vcc));
defparam a_valid.is_wysiwyg = "true";
defparam a_valid.power_up = "low";

fiftyfivenm_lcell_comb \Mux2~0 (
	.dataa(\in_ready_d1~q ),
	.datab(\state_d1[0]~q ),
	.datac(\state_register[0]~q ),
	.datad(\a_valid~q ),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'h1BE4;
defparam \Mux2~0 .sum_lutc_input = "datac";

dffeas \state_register[0] (
	.clk(clk),
	.d(\Mux2~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state_register[0]~q ),
	.prn(vcc));
defparam \state_register[0] .is_wysiwyg = "true";
defparam \state_register[0] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[0]~0 (
	.dataa(\a_data1[0]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[0]~0_combout ),
	.cout());
defparam \b_data[0]~0 .lut_mask = 16'h88A0;
defparam \b_data[0]~0 .sum_lutc_input = "datac";

dffeas \a_data1[1] (
	.clk(clk),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data1[1]~q ),
	.prn(vcc));
defparam \a_data1[1] .is_wysiwyg = "true";
defparam \a_data1[1] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[1]~1 (
	.dataa(\a_data1[1]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[1]~1_combout ),
	.cout());
defparam \b_data[1]~1 .lut_mask = 16'h88A0;
defparam \b_data[1]~1 .sum_lutc_input = "datac";

dffeas \a_data1[2] (
	.clk(clk),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data1[2]~q ),
	.prn(vcc));
defparam \a_data1[2] .is_wysiwyg = "true";
defparam \a_data1[2] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[2]~2 (
	.dataa(\a_data1[2]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[2]~2_combout ),
	.cout());
defparam \b_data[2]~2 .lut_mask = 16'h88A0;
defparam \b_data[2]~2 .sum_lutc_input = "datac";

dffeas \a_data1[3] (
	.clk(clk),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data1[3]~q ),
	.prn(vcc));
defparam \a_data1[3] .is_wysiwyg = "true";
defparam \a_data1[3] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[3]~3 (
	.dataa(\a_data1[3]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[3]~3_combout ),
	.cout());
defparam \b_data[3]~3 .lut_mask = 16'h88A0;
defparam \b_data[3]~3 .sum_lutc_input = "datac";

dffeas \a_data1[4] (
	.clk(clk),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data1[4]~q ),
	.prn(vcc));
defparam \a_data1[4] .is_wysiwyg = "true";
defparam \a_data1[4] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[4]~4 (
	.dataa(\a_data1[4]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[4]~4_combout ),
	.cout());
defparam \b_data[4]~4 .lut_mask = 16'h88A0;
defparam \b_data[4]~4 .sum_lutc_input = "datac";

dffeas \a_data1[5] (
	.clk(clk),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data1[5]~q ),
	.prn(vcc));
defparam \a_data1[5] .is_wysiwyg = "true";
defparam \a_data1[5] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[5]~5 (
	.dataa(\a_data1[5]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[5]~5_combout ),
	.cout());
defparam \b_data[5]~5 .lut_mask = 16'h88A0;
defparam \b_data[5]~5 .sum_lutc_input = "datac";

dffeas \a_data1[6] (
	.clk(clk),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data1[6]~q ),
	.prn(vcc));
defparam \a_data1[6] .is_wysiwyg = "true";
defparam \a_data1[6] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[6]~6 (
	.dataa(\a_data1[6]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[6]~6_combout ),
	.cout());
defparam \b_data[6]~6 .lut_mask = 16'h88A0;
defparam \b_data[6]~6 .sum_lutc_input = "datac";

dffeas \a_data1[7] (
	.clk(clk),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data1[7]~q ),
	.prn(vcc));
defparam \a_data1[7] .is_wysiwyg = "true";
defparam \a_data1[7] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[7]~7 (
	.dataa(\a_data1[7]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[7]~7_combout ),
	.cout());
defparam \b_data[7]~7 .lut_mask = 16'h88A0;
defparam \b_data[7]~7 .sum_lutc_input = "datac";

dffeas \a_data1[8] (
	.clk(clk),
	.d(in_data[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data1[8]~q ),
	.prn(vcc));
defparam \a_data1[8] .is_wysiwyg = "true";
defparam \a_data1[8] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[8]~8 (
	.dataa(\a_data1[8]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[8]~8_combout ),
	.cout());
defparam \b_data[8]~8 .lut_mask = 16'h88A0;
defparam \b_data[8]~8 .sum_lutc_input = "datac";

dffeas \a_data1[9] (
	.clk(clk),
	.d(in_data[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data1[9]~q ),
	.prn(vcc));
defparam \a_data1[9] .is_wysiwyg = "true";
defparam \a_data1[9] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[9]~9 (
	.dataa(\a_data1[9]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[9]~9_combout ),
	.cout());
defparam \b_data[9]~9 .lut_mask = 16'h88A0;
defparam \b_data[9]~9 .sum_lutc_input = "datac";

dffeas \a_data1[10] (
	.clk(clk),
	.d(in_data[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data1[10]~q ),
	.prn(vcc));
defparam \a_data1[10] .is_wysiwyg = "true";
defparam \a_data1[10] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[10]~10 (
	.dataa(\a_data1[10]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[10]~10_combout ),
	.cout());
defparam \b_data[10]~10 .lut_mask = 16'h88A0;
defparam \b_data[10]~10 .sum_lutc_input = "datac";

dffeas \a_data1[11] (
	.clk(clk),
	.d(in_data[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data1[11]~q ),
	.prn(vcc));
defparam \a_data1[11] .is_wysiwyg = "true";
defparam \a_data1[11] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[11]~11 (
	.dataa(\a_data1[11]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[11]~11_combout ),
	.cout());
defparam \b_data[11]~11 .lut_mask = 16'h88A0;
defparam \b_data[11]~11 .sum_lutc_input = "datac";

dffeas \a_data0[0] (
	.clk(clk),
	.d(in_data[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data0[0]~q ),
	.prn(vcc));
defparam \a_data0[0] .is_wysiwyg = "true";
defparam \a_data0[0] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[12]~12 (
	.dataa(\a_data0[0]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[12]~12_combout ),
	.cout());
defparam \b_data[12]~12 .lut_mask = 16'h88A0;
defparam \b_data[12]~12 .sum_lutc_input = "datac";

dffeas \a_data0[1] (
	.clk(clk),
	.d(in_data[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data0[1]~q ),
	.prn(vcc));
defparam \a_data0[1] .is_wysiwyg = "true";
defparam \a_data0[1] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[13]~13 (
	.dataa(\a_data0[1]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[13]~13_combout ),
	.cout());
defparam \b_data[13]~13 .lut_mask = 16'h88A0;
defparam \b_data[13]~13 .sum_lutc_input = "datac";

dffeas \a_data0[2] (
	.clk(clk),
	.d(in_data[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data0[2]~q ),
	.prn(vcc));
defparam \a_data0[2] .is_wysiwyg = "true";
defparam \a_data0[2] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[14]~14 (
	.dataa(\a_data0[2]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[14]~14_combout ),
	.cout());
defparam \b_data[14]~14 .lut_mask = 16'h88A0;
defparam \b_data[14]~14 .sum_lutc_input = "datac";

dffeas \a_data0[3] (
	.clk(clk),
	.d(in_data[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data0[3]~q ),
	.prn(vcc));
defparam \a_data0[3] .is_wysiwyg = "true";
defparam \a_data0[3] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[15]~15 (
	.dataa(\a_data0[3]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[15]~15_combout ),
	.cout());
defparam \b_data[15]~15 .lut_mask = 16'h88A0;
defparam \b_data[15]~15 .sum_lutc_input = "datac";

dffeas \a_data0[4] (
	.clk(clk),
	.d(in_data[16]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data0[4]~q ),
	.prn(vcc));
defparam \a_data0[4] .is_wysiwyg = "true";
defparam \a_data0[4] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[16]~16 (
	.dataa(\a_data0[4]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[16]~16_combout ),
	.cout());
defparam \b_data[16]~16 .lut_mask = 16'h88A0;
defparam \b_data[16]~16 .sum_lutc_input = "datac";

dffeas \a_data0[5] (
	.clk(clk),
	.d(in_data[17]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data0[5]~q ),
	.prn(vcc));
defparam \a_data0[5] .is_wysiwyg = "true";
defparam \a_data0[5] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[17]~17 (
	.dataa(\a_data0[5]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[17]~17_combout ),
	.cout());
defparam \b_data[17]~17 .lut_mask = 16'h88A0;
defparam \b_data[17]~17 .sum_lutc_input = "datac";

dffeas \a_data0[6] (
	.clk(clk),
	.d(in_data[18]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data0[6]~q ),
	.prn(vcc));
defparam \a_data0[6] .is_wysiwyg = "true";
defparam \a_data0[6] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[18]~18 (
	.dataa(\a_data0[6]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[18]~18_combout ),
	.cout());
defparam \b_data[18]~18 .lut_mask = 16'h88A0;
defparam \b_data[18]~18 .sum_lutc_input = "datac";

dffeas \a_data0[7] (
	.clk(clk),
	.d(in_data[19]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data0[7]~q ),
	.prn(vcc));
defparam \a_data0[7] .is_wysiwyg = "true";
defparam \a_data0[7] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[19]~19 (
	.dataa(\a_data0[7]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[19]~19_combout ),
	.cout());
defparam \b_data[19]~19 .lut_mask = 16'h88A0;
defparam \b_data[19]~19 .sum_lutc_input = "datac";

dffeas \a_data0[8] (
	.clk(clk),
	.d(in_data[20]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data0[8]~q ),
	.prn(vcc));
defparam \a_data0[8] .is_wysiwyg = "true";
defparam \a_data0[8] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[20]~20 (
	.dataa(\a_data0[8]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[20]~20_combout ),
	.cout());
defparam \b_data[20]~20 .lut_mask = 16'h88A0;
defparam \b_data[20]~20 .sum_lutc_input = "datac";

dffeas \a_data0[9] (
	.clk(clk),
	.d(in_data[21]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data0[9]~q ),
	.prn(vcc));
defparam \a_data0[9] .is_wysiwyg = "true";
defparam \a_data0[9] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[21]~21 (
	.dataa(\a_data0[9]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[21]~21_combout ),
	.cout());
defparam \b_data[21]~21 .lut_mask = 16'h88A0;
defparam \b_data[21]~21 .sum_lutc_input = "datac";

dffeas \a_data0[10] (
	.clk(clk),
	.d(in_data[22]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data0[10]~q ),
	.prn(vcc));
defparam \a_data0[10] .is_wysiwyg = "true";
defparam \a_data0[10] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[22]~22 (
	.dataa(\a_data0[10]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[22]~22_combout ),
	.cout());
defparam \b_data[22]~22 .lut_mask = 16'h88A0;
defparam \b_data[22]~22 .sum_lutc_input = "datac";

dffeas \a_data0[11] (
	.clk(clk),
	.d(in_data[23]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\a_data0[11]~q ),
	.prn(vcc));
defparam \a_data0[11] .is_wysiwyg = "true";
defparam \a_data0[11] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[23]~23 (
	.dataa(\a_data0[11]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[23]~23_combout ),
	.cout());
defparam \b_data[23]~23 .lut_mask = 16'h88A0;
defparam \b_data[23]~23 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux5~0 (
	.dataa(\a_valid~q ),
	.datab(\in_ready_d1~q ),
	.datac(\state_d1[0]~q ),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'h028A;
defparam \Mux5~0 .sum_lutc_input = "datac";

dffeas \data1_register[0] (
	.clk(clk),
	.d(\a_data1[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data1_register[0]~q ),
	.prn(vcc));
defparam \data1_register[0] .is_wysiwyg = "true";
defparam \data1_register[0] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[24]~24 (
	.dataa(\data1_register[0]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[24]~24_combout ),
	.cout());
defparam \b_data[24]~24 .lut_mask = 16'h88A0;
defparam \b_data[24]~24 .sum_lutc_input = "datac";

dffeas \data1_register[1] (
	.clk(clk),
	.d(\a_data1[1]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data1_register[1]~q ),
	.prn(vcc));
defparam \data1_register[1] .is_wysiwyg = "true";
defparam \data1_register[1] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[25]~25 (
	.dataa(\data1_register[1]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[25]~25_combout ),
	.cout());
defparam \b_data[25]~25 .lut_mask = 16'h88A0;
defparam \b_data[25]~25 .sum_lutc_input = "datac";

dffeas \data1_register[2] (
	.clk(clk),
	.d(\a_data1[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data1_register[2]~q ),
	.prn(vcc));
defparam \data1_register[2] .is_wysiwyg = "true";
defparam \data1_register[2] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[26]~26 (
	.dataa(\data1_register[2]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[26]~26_combout ),
	.cout());
defparam \b_data[26]~26 .lut_mask = 16'h88A0;
defparam \b_data[26]~26 .sum_lutc_input = "datac";

dffeas \data1_register[3] (
	.clk(clk),
	.d(\a_data1[3]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data1_register[3]~q ),
	.prn(vcc));
defparam \data1_register[3] .is_wysiwyg = "true";
defparam \data1_register[3] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[27]~27 (
	.dataa(\data1_register[3]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[27]~27_combout ),
	.cout());
defparam \b_data[27]~27 .lut_mask = 16'h88A0;
defparam \b_data[27]~27 .sum_lutc_input = "datac";

dffeas \data1_register[4] (
	.clk(clk),
	.d(\a_data1[4]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data1_register[4]~q ),
	.prn(vcc));
defparam \data1_register[4] .is_wysiwyg = "true";
defparam \data1_register[4] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[28]~28 (
	.dataa(\data1_register[4]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[28]~28_combout ),
	.cout());
defparam \b_data[28]~28 .lut_mask = 16'h88A0;
defparam \b_data[28]~28 .sum_lutc_input = "datac";

dffeas \data1_register[5] (
	.clk(clk),
	.d(\a_data1[5]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data1_register[5]~q ),
	.prn(vcc));
defparam \data1_register[5] .is_wysiwyg = "true";
defparam \data1_register[5] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[29]~29 (
	.dataa(\data1_register[5]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[29]~29_combout ),
	.cout());
defparam \b_data[29]~29 .lut_mask = 16'h88A0;
defparam \b_data[29]~29 .sum_lutc_input = "datac";

dffeas \data1_register[6] (
	.clk(clk),
	.d(\a_data1[6]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data1_register[6]~q ),
	.prn(vcc));
defparam \data1_register[6] .is_wysiwyg = "true";
defparam \data1_register[6] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[30]~30 (
	.dataa(\data1_register[6]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[30]~30_combout ),
	.cout());
defparam \b_data[30]~30 .lut_mask = 16'h88A0;
defparam \b_data[30]~30 .sum_lutc_input = "datac";

dffeas \data1_register[7] (
	.clk(clk),
	.d(\a_data1[7]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data1_register[7]~q ),
	.prn(vcc));
defparam \data1_register[7] .is_wysiwyg = "true";
defparam \data1_register[7] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[31]~31 (
	.dataa(\data1_register[7]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[31]~31_combout ),
	.cout());
defparam \b_data[31]~31 .lut_mask = 16'h88A0;
defparam \b_data[31]~31 .sum_lutc_input = "datac";

dffeas \data1_register[8] (
	.clk(clk),
	.d(\a_data1[8]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data1_register[8]~q ),
	.prn(vcc));
defparam \data1_register[8] .is_wysiwyg = "true";
defparam \data1_register[8] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[32]~32 (
	.dataa(\data1_register[8]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[32]~32_combout ),
	.cout());
defparam \b_data[32]~32 .lut_mask = 16'h88A0;
defparam \b_data[32]~32 .sum_lutc_input = "datac";

dffeas \data1_register[9] (
	.clk(clk),
	.d(\a_data1[9]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data1_register[9]~q ),
	.prn(vcc));
defparam \data1_register[9] .is_wysiwyg = "true";
defparam \data1_register[9] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[33]~33 (
	.dataa(\data1_register[9]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[33]~33_combout ),
	.cout());
defparam \b_data[33]~33 .lut_mask = 16'h88A0;
defparam \b_data[33]~33 .sum_lutc_input = "datac";

dffeas \data1_register[10] (
	.clk(clk),
	.d(\a_data1[10]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data1_register[10]~q ),
	.prn(vcc));
defparam \data1_register[10] .is_wysiwyg = "true";
defparam \data1_register[10] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[34]~34 (
	.dataa(\data1_register[10]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[34]~34_combout ),
	.cout());
defparam \b_data[34]~34 .lut_mask = 16'h88A0;
defparam \b_data[34]~34 .sum_lutc_input = "datac";

dffeas \data1_register[11] (
	.clk(clk),
	.d(\a_data1[11]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data1_register[11]~q ),
	.prn(vcc));
defparam \data1_register[11] .is_wysiwyg = "true";
defparam \data1_register[11] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[35]~35 (
	.dataa(\data1_register[11]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[35]~35_combout ),
	.cout());
defparam \b_data[35]~35 .lut_mask = 16'h88A0;
defparam \b_data[35]~35 .sum_lutc_input = "datac";

dffeas \data0_register[0] (
	.clk(clk),
	.d(\a_data0[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data0_register[0]~q ),
	.prn(vcc));
defparam \data0_register[0] .is_wysiwyg = "true";
defparam \data0_register[0] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[36]~36 (
	.dataa(\data0_register[0]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[36]~36_combout ),
	.cout());
defparam \b_data[36]~36 .lut_mask = 16'h88A0;
defparam \b_data[36]~36 .sum_lutc_input = "datac";

dffeas \data0_register[1] (
	.clk(clk),
	.d(\a_data0[1]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data0_register[1]~q ),
	.prn(vcc));
defparam \data0_register[1] .is_wysiwyg = "true";
defparam \data0_register[1] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[37]~37 (
	.dataa(\data0_register[1]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[37]~37_combout ),
	.cout());
defparam \b_data[37]~37 .lut_mask = 16'h88A0;
defparam \b_data[37]~37 .sum_lutc_input = "datac";

dffeas \data0_register[2] (
	.clk(clk),
	.d(\a_data0[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data0_register[2]~q ),
	.prn(vcc));
defparam \data0_register[2] .is_wysiwyg = "true";
defparam \data0_register[2] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[38]~38 (
	.dataa(\data0_register[2]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[38]~38_combout ),
	.cout());
defparam \b_data[38]~38 .lut_mask = 16'h88A0;
defparam \b_data[38]~38 .sum_lutc_input = "datac";

dffeas \data0_register[3] (
	.clk(clk),
	.d(\a_data0[3]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data0_register[3]~q ),
	.prn(vcc));
defparam \data0_register[3] .is_wysiwyg = "true";
defparam \data0_register[3] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[39]~39 (
	.dataa(\data0_register[3]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[39]~39_combout ),
	.cout());
defparam \b_data[39]~39 .lut_mask = 16'h88A0;
defparam \b_data[39]~39 .sum_lutc_input = "datac";

dffeas \data0_register[4] (
	.clk(clk),
	.d(\a_data0[4]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data0_register[4]~q ),
	.prn(vcc));
defparam \data0_register[4] .is_wysiwyg = "true";
defparam \data0_register[4] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[40]~40 (
	.dataa(\data0_register[4]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[40]~40_combout ),
	.cout());
defparam \b_data[40]~40 .lut_mask = 16'h88A0;
defparam \b_data[40]~40 .sum_lutc_input = "datac";

dffeas \data0_register[5] (
	.clk(clk),
	.d(\a_data0[5]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data0_register[5]~q ),
	.prn(vcc));
defparam \data0_register[5] .is_wysiwyg = "true";
defparam \data0_register[5] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[41]~41 (
	.dataa(\data0_register[5]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[41]~41_combout ),
	.cout());
defparam \b_data[41]~41 .lut_mask = 16'h88A0;
defparam \b_data[41]~41 .sum_lutc_input = "datac";

dffeas \data0_register[6] (
	.clk(clk),
	.d(\a_data0[6]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data0_register[6]~q ),
	.prn(vcc));
defparam \data0_register[6] .is_wysiwyg = "true";
defparam \data0_register[6] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[42]~42 (
	.dataa(\data0_register[6]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[42]~42_combout ),
	.cout());
defparam \b_data[42]~42 .lut_mask = 16'h88A0;
defparam \b_data[42]~42 .sum_lutc_input = "datac";

dffeas \data0_register[7] (
	.clk(clk),
	.d(\a_data0[7]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data0_register[7]~q ),
	.prn(vcc));
defparam \data0_register[7] .is_wysiwyg = "true";
defparam \data0_register[7] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[43]~43 (
	.dataa(\data0_register[7]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[43]~43_combout ),
	.cout());
defparam \b_data[43]~43 .lut_mask = 16'h88A0;
defparam \b_data[43]~43 .sum_lutc_input = "datac";

dffeas \data0_register[8] (
	.clk(clk),
	.d(\a_data0[8]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data0_register[8]~q ),
	.prn(vcc));
defparam \data0_register[8] .is_wysiwyg = "true";
defparam \data0_register[8] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[44]~44 (
	.dataa(\data0_register[8]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[44]~44_combout ),
	.cout());
defparam \b_data[44]~44 .lut_mask = 16'h88A0;
defparam \b_data[44]~44 .sum_lutc_input = "datac";

dffeas \data0_register[9] (
	.clk(clk),
	.d(\a_data0[9]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data0_register[9]~q ),
	.prn(vcc));
defparam \data0_register[9] .is_wysiwyg = "true";
defparam \data0_register[9] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[45]~45 (
	.dataa(\data0_register[9]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[45]~45_combout ),
	.cout());
defparam \b_data[45]~45 .lut_mask = 16'h88A0;
defparam \b_data[45]~45 .sum_lutc_input = "datac";

dffeas \data0_register[10] (
	.clk(clk),
	.d(\a_data0[10]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data0_register[10]~q ),
	.prn(vcc));
defparam \data0_register[10] .is_wysiwyg = "true";
defparam \data0_register[10] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[46]~46 (
	.dataa(\data0_register[10]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[46]~46_combout ),
	.cout());
defparam \b_data[46]~46 .lut_mask = 16'h88A0;
defparam \b_data[46]~46 .sum_lutc_input = "datac";

dffeas \data0_register[11] (
	.clk(clk),
	.d(\a_data0[11]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux5~0_combout ),
	.q(\data0_register[11]~q ),
	.prn(vcc));
defparam \data0_register[11] .is_wysiwyg = "true";
defparam \data0_register[11] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[47]~47 (
	.dataa(\data0_register[11]~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\b_data[47]~47_combout ),
	.cout());
defparam \b_data[47]~47 .lut_mask = 16'h88A0;
defparam \b_data[47]~47 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux3~0 (
	.dataa(\a_valid~q ),
	.datab(\state_register[0]~q ),
	.datac(\state_d1[0]~q ),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'h88A0;
defparam \Mux3~0 .sum_lutc_input = "datac";

endmodule

module lms_dsp_lms_dsp_avalon_st_adapter_001 (
	altera_reset_synchronizer_int_chain_out,
	out_valid,
	valid_reg,
	out_data_21,
	out_data_20,
	out_data_19,
	out_data_18,
	out_data_17,
	out_data_16,
	out_data_15,
	out_data_14,
	out_data_12,
	out_data_13,
	out_data_9,
	out_data_8,
	out_data_7,
	out_data_6,
	out_data_5,
	out_data_4,
	out_data_3,
	out_data_2,
	out_data_0,
	out_data_1,
	out_data_11,
	out_data_10,
	out_data_23,
	out_data_22,
	data_reg_21,
	data_reg_45,
	data_reg_20,
	data_reg_44,
	data_reg_19,
	data_reg_43,
	data_reg_18,
	data_reg_42,
	data_reg_17,
	data_reg_41,
	data_reg_16,
	data_reg_40,
	data_reg_15,
	data_reg_39,
	data_reg_14,
	data_reg_38,
	data_reg_12,
	data_reg_36,
	data_reg_13,
	data_reg_37,
	data_reg_9,
	data_reg_33,
	data_reg_8,
	data_reg_32,
	data_reg_7,
	data_reg_31,
	data_reg_6,
	data_reg_30,
	data_reg_5,
	data_reg_29,
	data_reg_4,
	data_reg_28,
	data_reg_3,
	data_reg_27,
	data_reg_2,
	data_reg_26,
	data_reg_0,
	data_reg_24,
	data_reg_1,
	data_reg_25,
	data_reg_11,
	data_reg_35,
	data_reg_10,
	data_reg_34,
	data_reg_23,
	data_reg_47,
	data_reg_22,
	data_reg_46,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	altera_reset_synchronizer_int_chain_out;
output 	out_valid;
input 	valid_reg;
output 	out_data_21;
output 	out_data_20;
output 	out_data_19;
output 	out_data_18;
output 	out_data_17;
output 	out_data_16;
output 	out_data_15;
output 	out_data_14;
output 	out_data_12;
output 	out_data_13;
output 	out_data_9;
output 	out_data_8;
output 	out_data_7;
output 	out_data_6;
output 	out_data_5;
output 	out_data_4;
output 	out_data_3;
output 	out_data_2;
output 	out_data_0;
output 	out_data_1;
output 	out_data_11;
output 	out_data_10;
output 	out_data_23;
output 	out_data_22;
input 	data_reg_21;
input 	data_reg_45;
input 	data_reg_20;
input 	data_reg_44;
input 	data_reg_19;
input 	data_reg_43;
input 	data_reg_18;
input 	data_reg_42;
input 	data_reg_17;
input 	data_reg_41;
input 	data_reg_16;
input 	data_reg_40;
input 	data_reg_15;
input 	data_reg_39;
input 	data_reg_14;
input 	data_reg_38;
input 	data_reg_12;
input 	data_reg_36;
input 	data_reg_13;
input 	data_reg_37;
input 	data_reg_9;
input 	data_reg_33;
input 	data_reg_8;
input 	data_reg_32;
input 	data_reg_7;
input 	data_reg_31;
input 	data_reg_6;
input 	data_reg_30;
input 	data_reg_5;
input 	data_reg_29;
input 	data_reg_4;
input 	data_reg_28;
input 	data_reg_3;
input 	data_reg_27;
input 	data_reg_2;
input 	data_reg_26;
input 	data_reg_0;
input 	data_reg_24;
input 	data_reg_1;
input 	data_reg_25;
input 	data_reg_11;
input 	data_reg_35;
input 	data_reg_10;
input 	data_reg_34;
input 	data_reg_23;
input 	data_reg_47;
input 	data_reg_22;
input 	data_reg_46;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



lms_dsp_lms_dsp_avalon_st_adapter_001_data_format_adapter_0 data_format_adapter_0(
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.out_valid1(out_valid),
	.in_valid(valid_reg),
	.out_data_21(out_data_21),
	.out_data_20(out_data_20),
	.out_data_19(out_data_19),
	.out_data_18(out_data_18),
	.out_data_17(out_data_17),
	.out_data_16(out_data_16),
	.out_data_15(out_data_15),
	.out_data_14(out_data_14),
	.out_data_12(out_data_12),
	.out_data_13(out_data_13),
	.out_data_9(out_data_9),
	.out_data_8(out_data_8),
	.out_data_7(out_data_7),
	.out_data_6(out_data_6),
	.out_data_5(out_data_5),
	.out_data_4(out_data_4),
	.out_data_3(out_data_3),
	.out_data_2(out_data_2),
	.out_data_0(out_data_0),
	.out_data_1(out_data_1),
	.out_data_11(out_data_11),
	.out_data_10(out_data_10),
	.out_data_23(out_data_23),
	.out_data_22(out_data_22),
	.in_data({data_reg_47,data_reg_46,data_reg_45,data_reg_44,data_reg_43,data_reg_42,data_reg_41,data_reg_40,data_reg_39,data_reg_38,data_reg_37,data_reg_36,data_reg_35,data_reg_34,data_reg_33,data_reg_32,data_reg_31,data_reg_30,data_reg_29,data_reg_28,data_reg_27,data_reg_26,data_reg_25,
data_reg_24,data_reg_23,data_reg_22,data_reg_21,data_reg_20,data_reg_19,data_reg_18,data_reg_17,data_reg_16,data_reg_15,data_reg_14,data_reg_13,data_reg_12,data_reg_11,data_reg_10,data_reg_9,data_reg_8,data_reg_7,data_reg_6,data_reg_5,data_reg_4,data_reg_3,data_reg_2,data_reg_1,
data_reg_0}),
	.clk(clk_clk));

endmodule

module lms_dsp_lms_dsp_avalon_st_adapter_001_data_format_adapter_0 (
	reset_n,
	out_valid1,
	in_valid,
	out_data_21,
	out_data_20,
	out_data_19,
	out_data_18,
	out_data_17,
	out_data_16,
	out_data_15,
	out_data_14,
	out_data_12,
	out_data_13,
	out_data_9,
	out_data_8,
	out_data_7,
	out_data_6,
	out_data_5,
	out_data_4,
	out_data_3,
	out_data_2,
	out_data_0,
	out_data_1,
	out_data_11,
	out_data_10,
	out_data_23,
	out_data_22,
	in_data,
	clk)/* synthesis synthesis_greybox=0 */;
input 	reset_n;
output 	out_valid1;
input 	in_valid;
output 	out_data_21;
output 	out_data_20;
output 	out_data_19;
output 	out_data_18;
output 	out_data_17;
output 	out_data_16;
output 	out_data_15;
output 	out_data_14;
output 	out_data_12;
output 	out_data_13;
output 	out_data_9;
output 	out_data_8;
output 	out_data_7;
output 	out_data_6;
output 	out_data_5;
output 	out_data_4;
output 	out_data_3;
output 	out_data_2;
output 	out_data_0;
output 	out_data_1;
output 	out_data_11;
output 	out_data_10;
output 	out_data_23;
output 	out_data_22;
input 	[47:0] in_data;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \state_register[0]~0_combout ;
wire \state_register[0]~q ;
wire \in_ready~combout ;
wire \a_valid~q ;
wire \a_data2[9]~q ;
wire \a_data0[9]~q ;
wire \b_data[21]~0_combout ;
wire \a_data2[8]~q ;
wire \a_data0[8]~q ;
wire \b_data[20]~1_combout ;
wire \a_data2[7]~q ;
wire \a_data0[7]~q ;
wire \b_data[19]~2_combout ;
wire \a_data2[6]~q ;
wire \a_data0[6]~q ;
wire \b_data[18]~3_combout ;
wire \a_data2[5]~q ;
wire \a_data0[5]~q ;
wire \b_data[17]~4_combout ;
wire \a_data2[4]~q ;
wire \a_data0[4]~q ;
wire \b_data[16]~5_combout ;
wire \a_data2[3]~q ;
wire \a_data0[3]~q ;
wire \b_data[15]~6_combout ;
wire \a_data2[2]~q ;
wire \a_data0[2]~q ;
wire \b_data[14]~7_combout ;
wire \a_data2[0]~q ;
wire \a_data0[0]~q ;
wire \b_data[12]~8_combout ;
wire \a_data2[1]~q ;
wire \a_data0[1]~q ;
wire \b_data[13]~9_combout ;
wire \a_data3[9]~q ;
wire \a_data1[9]~q ;
wire \b_data[9]~10_combout ;
wire \a_data3[8]~q ;
wire \a_data1[8]~q ;
wire \b_data[8]~11_combout ;
wire \a_data3[7]~q ;
wire \a_data1[7]~q ;
wire \b_data[7]~12_combout ;
wire \a_data3[6]~q ;
wire \a_data1[6]~q ;
wire \b_data[6]~13_combout ;
wire \a_data3[5]~q ;
wire \a_data1[5]~q ;
wire \b_data[5]~14_combout ;
wire \a_data3[4]~q ;
wire \a_data1[4]~q ;
wire \b_data[4]~15_combout ;
wire \a_data3[3]~q ;
wire \a_data1[3]~q ;
wire \b_data[3]~16_combout ;
wire \a_data3[2]~q ;
wire \a_data1[2]~q ;
wire \b_data[2]~17_combout ;
wire \a_data3[0]~q ;
wire \a_data1[0]~q ;
wire \b_data[0]~18_combout ;
wire \a_data3[1]~q ;
wire \a_data1[1]~q ;
wire \b_data[1]~19_combout ;
wire \a_data3[11]~q ;
wire \a_data1[11]~q ;
wire \b_data[11]~20_combout ;
wire \a_data3[10]~q ;
wire \a_data1[10]~q ;
wire \b_data[10]~21_combout ;
wire \a_data2[11]~q ;
wire \a_data0[11]~q ;
wire \b_data[23]~22_combout ;
wire \a_data2[10]~q ;
wire \a_data0[10]~q ;
wire \b_data[22]~23_combout ;


dffeas out_valid(
	.clk(clk),
	.d(\a_valid~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

dffeas \out_data[21] (
	.clk(clk),
	.d(\b_data[21]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_21),
	.prn(vcc));
defparam \out_data[21] .is_wysiwyg = "true";
defparam \out_data[21] .power_up = "low";

dffeas \out_data[20] (
	.clk(clk),
	.d(\b_data[20]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_20),
	.prn(vcc));
defparam \out_data[20] .is_wysiwyg = "true";
defparam \out_data[20] .power_up = "low";

dffeas \out_data[19] (
	.clk(clk),
	.d(\b_data[19]~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_19),
	.prn(vcc));
defparam \out_data[19] .is_wysiwyg = "true";
defparam \out_data[19] .power_up = "low";

dffeas \out_data[18] (
	.clk(clk),
	.d(\b_data[18]~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_18),
	.prn(vcc));
defparam \out_data[18] .is_wysiwyg = "true";
defparam \out_data[18] .power_up = "low";

dffeas \out_data[17] (
	.clk(clk),
	.d(\b_data[17]~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_17),
	.prn(vcc));
defparam \out_data[17] .is_wysiwyg = "true";
defparam \out_data[17] .power_up = "low";

dffeas \out_data[16] (
	.clk(clk),
	.d(\b_data[16]~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_16),
	.prn(vcc));
defparam \out_data[16] .is_wysiwyg = "true";
defparam \out_data[16] .power_up = "low";

dffeas \out_data[15] (
	.clk(clk),
	.d(\b_data[15]~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_15),
	.prn(vcc));
defparam \out_data[15] .is_wysiwyg = "true";
defparam \out_data[15] .power_up = "low";

dffeas \out_data[14] (
	.clk(clk),
	.d(\b_data[14]~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_14),
	.prn(vcc));
defparam \out_data[14] .is_wysiwyg = "true";
defparam \out_data[14] .power_up = "low";

dffeas \out_data[12] (
	.clk(clk),
	.d(\b_data[12]~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_12),
	.prn(vcc));
defparam \out_data[12] .is_wysiwyg = "true";
defparam \out_data[12] .power_up = "low";

dffeas \out_data[13] (
	.clk(clk),
	.d(\b_data[13]~9_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_13),
	.prn(vcc));
defparam \out_data[13] .is_wysiwyg = "true";
defparam \out_data[13] .power_up = "low";

dffeas \out_data[9] (
	.clk(clk),
	.d(\b_data[9]~10_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_9),
	.prn(vcc));
defparam \out_data[9] .is_wysiwyg = "true";
defparam \out_data[9] .power_up = "low";

dffeas \out_data[8] (
	.clk(clk),
	.d(\b_data[8]~11_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_8),
	.prn(vcc));
defparam \out_data[8] .is_wysiwyg = "true";
defparam \out_data[8] .power_up = "low";

dffeas \out_data[7] (
	.clk(clk),
	.d(\b_data[7]~12_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_7),
	.prn(vcc));
defparam \out_data[7] .is_wysiwyg = "true";
defparam \out_data[7] .power_up = "low";

dffeas \out_data[6] (
	.clk(clk),
	.d(\b_data[6]~13_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_6),
	.prn(vcc));
defparam \out_data[6] .is_wysiwyg = "true";
defparam \out_data[6] .power_up = "low";

dffeas \out_data[5] (
	.clk(clk),
	.d(\b_data[5]~14_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_5),
	.prn(vcc));
defparam \out_data[5] .is_wysiwyg = "true";
defparam \out_data[5] .power_up = "low";

dffeas \out_data[4] (
	.clk(clk),
	.d(\b_data[4]~15_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_4),
	.prn(vcc));
defparam \out_data[4] .is_wysiwyg = "true";
defparam \out_data[4] .power_up = "low";

dffeas \out_data[3] (
	.clk(clk),
	.d(\b_data[3]~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_3),
	.prn(vcc));
defparam \out_data[3] .is_wysiwyg = "true";
defparam \out_data[3] .power_up = "low";

dffeas \out_data[2] (
	.clk(clk),
	.d(\b_data[2]~17_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_2),
	.prn(vcc));
defparam \out_data[2] .is_wysiwyg = "true";
defparam \out_data[2] .power_up = "low";

dffeas \out_data[0] (
	.clk(clk),
	.d(\b_data[0]~18_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_0),
	.prn(vcc));
defparam \out_data[0] .is_wysiwyg = "true";
defparam \out_data[0] .power_up = "low";

dffeas \out_data[1] (
	.clk(clk),
	.d(\b_data[1]~19_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_1),
	.prn(vcc));
defparam \out_data[1] .is_wysiwyg = "true";
defparam \out_data[1] .power_up = "low";

dffeas \out_data[11] (
	.clk(clk),
	.d(\b_data[11]~20_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_11),
	.prn(vcc));
defparam \out_data[11] .is_wysiwyg = "true";
defparam \out_data[11] .power_up = "low";

dffeas \out_data[10] (
	.clk(clk),
	.d(\b_data[10]~21_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_10),
	.prn(vcc));
defparam \out_data[10] .is_wysiwyg = "true";
defparam \out_data[10] .power_up = "low";

dffeas \out_data[23] (
	.clk(clk),
	.d(\b_data[23]~22_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_23),
	.prn(vcc));
defparam \out_data[23] .is_wysiwyg = "true";
defparam \out_data[23] .power_up = "low";

dffeas \out_data[22] (
	.clk(clk),
	.d(\b_data[22]~23_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_22),
	.prn(vcc));
defparam \out_data[22] .is_wysiwyg = "true";
defparam \out_data[22] .power_up = "low";

fiftyfivenm_lcell_comb \state_register[0]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\a_valid~q ),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\state_register[0]~0_combout ),
	.cout());
defparam \state_register[0]~0 .lut_mask = 16'h0FF0;
defparam \state_register[0]~0 .sum_lutc_input = "datac";

dffeas \state_register[0] (
	.clk(clk),
	.d(\state_register[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state_register[0]~q ),
	.prn(vcc));
defparam \state_register[0] .is_wysiwyg = "true";
defparam \state_register[0] .power_up = "low";

fiftyfivenm_lcell_comb in_ready(
	.dataa(\state_register[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\a_valid~q ),
	.cin(gnd),
	.combout(\in_ready~combout ),
	.cout());
defparam in_ready.lut_mask = 16'hAAFF;
defparam in_ready.sum_lutc_input = "datac";

dffeas a_valid(
	.clk(clk),
	.d(in_valid),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_valid~q ),
	.prn(vcc));
defparam a_valid.is_wysiwyg = "true";
defparam a_valid.power_up = "low";

dffeas \a_data2[9] (
	.clk(clk),
	.d(in_data[21]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data2[9]~q ),
	.prn(vcc));
defparam \a_data2[9] .is_wysiwyg = "true";
defparam \a_data2[9] .power_up = "low";

dffeas \a_data0[9] (
	.clk(clk),
	.d(in_data[45]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data0[9]~q ),
	.prn(vcc));
defparam \a_data0[9] .is_wysiwyg = "true";
defparam \a_data0[9] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[21]~0 (
	.dataa(\a_data2[9]~q ),
	.datab(\a_data0[9]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[21]~0_combout ),
	.cout());
defparam \b_data[21]~0 .lut_mask = 16'hAACC;
defparam \b_data[21]~0 .sum_lutc_input = "datac";

dffeas \a_data2[8] (
	.clk(clk),
	.d(in_data[20]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data2[8]~q ),
	.prn(vcc));
defparam \a_data2[8] .is_wysiwyg = "true";
defparam \a_data2[8] .power_up = "low";

dffeas \a_data0[8] (
	.clk(clk),
	.d(in_data[44]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data0[8]~q ),
	.prn(vcc));
defparam \a_data0[8] .is_wysiwyg = "true";
defparam \a_data0[8] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[20]~1 (
	.dataa(\a_data2[8]~q ),
	.datab(\a_data0[8]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[20]~1_combout ),
	.cout());
defparam \b_data[20]~1 .lut_mask = 16'hAACC;
defparam \b_data[20]~1 .sum_lutc_input = "datac";

dffeas \a_data2[7] (
	.clk(clk),
	.d(in_data[19]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data2[7]~q ),
	.prn(vcc));
defparam \a_data2[7] .is_wysiwyg = "true";
defparam \a_data2[7] .power_up = "low";

dffeas \a_data0[7] (
	.clk(clk),
	.d(in_data[43]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data0[7]~q ),
	.prn(vcc));
defparam \a_data0[7] .is_wysiwyg = "true";
defparam \a_data0[7] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[19]~2 (
	.dataa(\a_data2[7]~q ),
	.datab(\a_data0[7]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[19]~2_combout ),
	.cout());
defparam \b_data[19]~2 .lut_mask = 16'hAACC;
defparam \b_data[19]~2 .sum_lutc_input = "datac";

dffeas \a_data2[6] (
	.clk(clk),
	.d(in_data[18]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data2[6]~q ),
	.prn(vcc));
defparam \a_data2[6] .is_wysiwyg = "true";
defparam \a_data2[6] .power_up = "low";

dffeas \a_data0[6] (
	.clk(clk),
	.d(in_data[42]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data0[6]~q ),
	.prn(vcc));
defparam \a_data0[6] .is_wysiwyg = "true";
defparam \a_data0[6] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[18]~3 (
	.dataa(\a_data2[6]~q ),
	.datab(\a_data0[6]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[18]~3_combout ),
	.cout());
defparam \b_data[18]~3 .lut_mask = 16'hAACC;
defparam \b_data[18]~3 .sum_lutc_input = "datac";

dffeas \a_data2[5] (
	.clk(clk),
	.d(in_data[17]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data2[5]~q ),
	.prn(vcc));
defparam \a_data2[5] .is_wysiwyg = "true";
defparam \a_data2[5] .power_up = "low";

dffeas \a_data0[5] (
	.clk(clk),
	.d(in_data[41]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data0[5]~q ),
	.prn(vcc));
defparam \a_data0[5] .is_wysiwyg = "true";
defparam \a_data0[5] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[17]~4 (
	.dataa(\a_data2[5]~q ),
	.datab(\a_data0[5]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[17]~4_combout ),
	.cout());
defparam \b_data[17]~4 .lut_mask = 16'hAACC;
defparam \b_data[17]~4 .sum_lutc_input = "datac";

dffeas \a_data2[4] (
	.clk(clk),
	.d(in_data[16]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data2[4]~q ),
	.prn(vcc));
defparam \a_data2[4] .is_wysiwyg = "true";
defparam \a_data2[4] .power_up = "low";

dffeas \a_data0[4] (
	.clk(clk),
	.d(in_data[40]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data0[4]~q ),
	.prn(vcc));
defparam \a_data0[4] .is_wysiwyg = "true";
defparam \a_data0[4] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[16]~5 (
	.dataa(\a_data2[4]~q ),
	.datab(\a_data0[4]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[16]~5_combout ),
	.cout());
defparam \b_data[16]~5 .lut_mask = 16'hAACC;
defparam \b_data[16]~5 .sum_lutc_input = "datac";

dffeas \a_data2[3] (
	.clk(clk),
	.d(in_data[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data2[3]~q ),
	.prn(vcc));
defparam \a_data2[3] .is_wysiwyg = "true";
defparam \a_data2[3] .power_up = "low";

dffeas \a_data0[3] (
	.clk(clk),
	.d(in_data[39]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data0[3]~q ),
	.prn(vcc));
defparam \a_data0[3] .is_wysiwyg = "true";
defparam \a_data0[3] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[15]~6 (
	.dataa(\a_data2[3]~q ),
	.datab(\a_data0[3]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[15]~6_combout ),
	.cout());
defparam \b_data[15]~6 .lut_mask = 16'hAACC;
defparam \b_data[15]~6 .sum_lutc_input = "datac";

dffeas \a_data2[2] (
	.clk(clk),
	.d(in_data[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data2[2]~q ),
	.prn(vcc));
defparam \a_data2[2] .is_wysiwyg = "true";
defparam \a_data2[2] .power_up = "low";

dffeas \a_data0[2] (
	.clk(clk),
	.d(in_data[38]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data0[2]~q ),
	.prn(vcc));
defparam \a_data0[2] .is_wysiwyg = "true";
defparam \a_data0[2] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[14]~7 (
	.dataa(\a_data2[2]~q ),
	.datab(\a_data0[2]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[14]~7_combout ),
	.cout());
defparam \b_data[14]~7 .lut_mask = 16'hAACC;
defparam \b_data[14]~7 .sum_lutc_input = "datac";

dffeas \a_data2[0] (
	.clk(clk),
	.d(in_data[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data2[0]~q ),
	.prn(vcc));
defparam \a_data2[0] .is_wysiwyg = "true";
defparam \a_data2[0] .power_up = "low";

dffeas \a_data0[0] (
	.clk(clk),
	.d(in_data[36]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data0[0]~q ),
	.prn(vcc));
defparam \a_data0[0] .is_wysiwyg = "true";
defparam \a_data0[0] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[12]~8 (
	.dataa(\a_data2[0]~q ),
	.datab(\a_data0[0]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[12]~8_combout ),
	.cout());
defparam \b_data[12]~8 .lut_mask = 16'hAACC;
defparam \b_data[12]~8 .sum_lutc_input = "datac";

dffeas \a_data2[1] (
	.clk(clk),
	.d(in_data[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data2[1]~q ),
	.prn(vcc));
defparam \a_data2[1] .is_wysiwyg = "true";
defparam \a_data2[1] .power_up = "low";

dffeas \a_data0[1] (
	.clk(clk),
	.d(in_data[37]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data0[1]~q ),
	.prn(vcc));
defparam \a_data0[1] .is_wysiwyg = "true";
defparam \a_data0[1] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[13]~9 (
	.dataa(\a_data2[1]~q ),
	.datab(\a_data0[1]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[13]~9_combout ),
	.cout());
defparam \b_data[13]~9 .lut_mask = 16'hAACC;
defparam \b_data[13]~9 .sum_lutc_input = "datac";

dffeas \a_data3[9] (
	.clk(clk),
	.d(in_data[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data3[9]~q ),
	.prn(vcc));
defparam \a_data3[9] .is_wysiwyg = "true";
defparam \a_data3[9] .power_up = "low";

dffeas \a_data1[9] (
	.clk(clk),
	.d(in_data[33]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data1[9]~q ),
	.prn(vcc));
defparam \a_data1[9] .is_wysiwyg = "true";
defparam \a_data1[9] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[9]~10 (
	.dataa(\a_data3[9]~q ),
	.datab(\a_data1[9]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[9]~10_combout ),
	.cout());
defparam \b_data[9]~10 .lut_mask = 16'hAACC;
defparam \b_data[9]~10 .sum_lutc_input = "datac";

dffeas \a_data3[8] (
	.clk(clk),
	.d(in_data[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data3[8]~q ),
	.prn(vcc));
defparam \a_data3[8] .is_wysiwyg = "true";
defparam \a_data3[8] .power_up = "low";

dffeas \a_data1[8] (
	.clk(clk),
	.d(in_data[32]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data1[8]~q ),
	.prn(vcc));
defparam \a_data1[8] .is_wysiwyg = "true";
defparam \a_data1[8] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[8]~11 (
	.dataa(\a_data3[8]~q ),
	.datab(\a_data1[8]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[8]~11_combout ),
	.cout());
defparam \b_data[8]~11 .lut_mask = 16'hAACC;
defparam \b_data[8]~11 .sum_lutc_input = "datac";

dffeas \a_data3[7] (
	.clk(clk),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data3[7]~q ),
	.prn(vcc));
defparam \a_data3[7] .is_wysiwyg = "true";
defparam \a_data3[7] .power_up = "low";

dffeas \a_data1[7] (
	.clk(clk),
	.d(in_data[31]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data1[7]~q ),
	.prn(vcc));
defparam \a_data1[7] .is_wysiwyg = "true";
defparam \a_data1[7] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[7]~12 (
	.dataa(\a_data3[7]~q ),
	.datab(\a_data1[7]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[7]~12_combout ),
	.cout());
defparam \b_data[7]~12 .lut_mask = 16'hAACC;
defparam \b_data[7]~12 .sum_lutc_input = "datac";

dffeas \a_data3[6] (
	.clk(clk),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data3[6]~q ),
	.prn(vcc));
defparam \a_data3[6] .is_wysiwyg = "true";
defparam \a_data3[6] .power_up = "low";

dffeas \a_data1[6] (
	.clk(clk),
	.d(in_data[30]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data1[6]~q ),
	.prn(vcc));
defparam \a_data1[6] .is_wysiwyg = "true";
defparam \a_data1[6] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[6]~13 (
	.dataa(\a_data3[6]~q ),
	.datab(\a_data1[6]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[6]~13_combout ),
	.cout());
defparam \b_data[6]~13 .lut_mask = 16'hAACC;
defparam \b_data[6]~13 .sum_lutc_input = "datac";

dffeas \a_data3[5] (
	.clk(clk),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data3[5]~q ),
	.prn(vcc));
defparam \a_data3[5] .is_wysiwyg = "true";
defparam \a_data3[5] .power_up = "low";

dffeas \a_data1[5] (
	.clk(clk),
	.d(in_data[29]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data1[5]~q ),
	.prn(vcc));
defparam \a_data1[5] .is_wysiwyg = "true";
defparam \a_data1[5] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[5]~14 (
	.dataa(\a_data3[5]~q ),
	.datab(\a_data1[5]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[5]~14_combout ),
	.cout());
defparam \b_data[5]~14 .lut_mask = 16'hAACC;
defparam \b_data[5]~14 .sum_lutc_input = "datac";

dffeas \a_data3[4] (
	.clk(clk),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data3[4]~q ),
	.prn(vcc));
defparam \a_data3[4] .is_wysiwyg = "true";
defparam \a_data3[4] .power_up = "low";

dffeas \a_data1[4] (
	.clk(clk),
	.d(in_data[28]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data1[4]~q ),
	.prn(vcc));
defparam \a_data1[4] .is_wysiwyg = "true";
defparam \a_data1[4] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[4]~15 (
	.dataa(\a_data3[4]~q ),
	.datab(\a_data1[4]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[4]~15_combout ),
	.cout());
defparam \b_data[4]~15 .lut_mask = 16'hAACC;
defparam \b_data[4]~15 .sum_lutc_input = "datac";

dffeas \a_data3[3] (
	.clk(clk),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data3[3]~q ),
	.prn(vcc));
defparam \a_data3[3] .is_wysiwyg = "true";
defparam \a_data3[3] .power_up = "low";

dffeas \a_data1[3] (
	.clk(clk),
	.d(in_data[27]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data1[3]~q ),
	.prn(vcc));
defparam \a_data1[3] .is_wysiwyg = "true";
defparam \a_data1[3] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[3]~16 (
	.dataa(\a_data3[3]~q ),
	.datab(\a_data1[3]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[3]~16_combout ),
	.cout());
defparam \b_data[3]~16 .lut_mask = 16'hAACC;
defparam \b_data[3]~16 .sum_lutc_input = "datac";

dffeas \a_data3[2] (
	.clk(clk),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data3[2]~q ),
	.prn(vcc));
defparam \a_data3[2] .is_wysiwyg = "true";
defparam \a_data3[2] .power_up = "low";

dffeas \a_data1[2] (
	.clk(clk),
	.d(in_data[26]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data1[2]~q ),
	.prn(vcc));
defparam \a_data1[2] .is_wysiwyg = "true";
defparam \a_data1[2] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[2]~17 (
	.dataa(\a_data3[2]~q ),
	.datab(\a_data1[2]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[2]~17_combout ),
	.cout());
defparam \b_data[2]~17 .lut_mask = 16'hAACC;
defparam \b_data[2]~17 .sum_lutc_input = "datac";

dffeas \a_data3[0] (
	.clk(clk),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data3[0]~q ),
	.prn(vcc));
defparam \a_data3[0] .is_wysiwyg = "true";
defparam \a_data3[0] .power_up = "low";

dffeas \a_data1[0] (
	.clk(clk),
	.d(in_data[24]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data1[0]~q ),
	.prn(vcc));
defparam \a_data1[0] .is_wysiwyg = "true";
defparam \a_data1[0] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[0]~18 (
	.dataa(\a_data3[0]~q ),
	.datab(\a_data1[0]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[0]~18_combout ),
	.cout());
defparam \b_data[0]~18 .lut_mask = 16'hAACC;
defparam \b_data[0]~18 .sum_lutc_input = "datac";

dffeas \a_data3[1] (
	.clk(clk),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data3[1]~q ),
	.prn(vcc));
defparam \a_data3[1] .is_wysiwyg = "true";
defparam \a_data3[1] .power_up = "low";

dffeas \a_data1[1] (
	.clk(clk),
	.d(in_data[25]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data1[1]~q ),
	.prn(vcc));
defparam \a_data1[1] .is_wysiwyg = "true";
defparam \a_data1[1] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[1]~19 (
	.dataa(\a_data3[1]~q ),
	.datab(\a_data1[1]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[1]~19_combout ),
	.cout());
defparam \b_data[1]~19 .lut_mask = 16'hAACC;
defparam \b_data[1]~19 .sum_lutc_input = "datac";

dffeas \a_data3[11] (
	.clk(clk),
	.d(in_data[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data3[11]~q ),
	.prn(vcc));
defparam \a_data3[11] .is_wysiwyg = "true";
defparam \a_data3[11] .power_up = "low";

dffeas \a_data1[11] (
	.clk(clk),
	.d(in_data[35]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data1[11]~q ),
	.prn(vcc));
defparam \a_data1[11] .is_wysiwyg = "true";
defparam \a_data1[11] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[11]~20 (
	.dataa(\a_data3[11]~q ),
	.datab(\a_data1[11]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[11]~20_combout ),
	.cout());
defparam \b_data[11]~20 .lut_mask = 16'hAACC;
defparam \b_data[11]~20 .sum_lutc_input = "datac";

dffeas \a_data3[10] (
	.clk(clk),
	.d(in_data[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data3[10]~q ),
	.prn(vcc));
defparam \a_data3[10] .is_wysiwyg = "true";
defparam \a_data3[10] .power_up = "low";

dffeas \a_data1[10] (
	.clk(clk),
	.d(in_data[34]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data1[10]~q ),
	.prn(vcc));
defparam \a_data1[10] .is_wysiwyg = "true";
defparam \a_data1[10] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[10]~21 (
	.dataa(\a_data3[10]~q ),
	.datab(\a_data1[10]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[10]~21_combout ),
	.cout());
defparam \b_data[10]~21 .lut_mask = 16'hAACC;
defparam \b_data[10]~21 .sum_lutc_input = "datac";

dffeas \a_data2[11] (
	.clk(clk),
	.d(in_data[23]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data2[11]~q ),
	.prn(vcc));
defparam \a_data2[11] .is_wysiwyg = "true";
defparam \a_data2[11] .power_up = "low";

dffeas \a_data0[11] (
	.clk(clk),
	.d(in_data[47]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data0[11]~q ),
	.prn(vcc));
defparam \a_data0[11] .is_wysiwyg = "true";
defparam \a_data0[11] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[23]~22 (
	.dataa(\a_data2[11]~q ),
	.datab(\a_data0[11]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[23]~22_combout ),
	.cout());
defparam \b_data[23]~22 .lut_mask = 16'hAACC;
defparam \b_data[23]~22 .sum_lutc_input = "datac";

dffeas \a_data2[10] (
	.clk(clk),
	.d(in_data[22]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data2[10]~q ),
	.prn(vcc));
defparam \a_data2[10] .is_wysiwyg = "true";
defparam \a_data2[10] .power_up = "low";

dffeas \a_data0[10] (
	.clk(clk),
	.d(in_data[46]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~combout ),
	.q(\a_data0[10]~q ),
	.prn(vcc));
defparam \a_data0[10] .is_wysiwyg = "true";
defparam \a_data0[10] .power_up = "low";

fiftyfivenm_lcell_comb \b_data[22]~23 (
	.dataa(\a_data2[10]~q ),
	.datab(\a_data0[10]~q ),
	.datac(gnd),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\b_data[22]~23_combout ),
	.cout());
defparam \b_data[22]~23 .lut_mask = 16'hAACC;
defparam \b_data[22]~23 .sum_lutc_input = "datac";

endmodule

module lms_dsp_lms_dsp_fir_compiler_ii_0 (
	reset_n,
	data_out_12,
	data_out_0,
	data_out_11,
	data_out_10,
	data_out_9,
	data_out_8,
	data_out_7,
	data_out_6,
	data_out_5,
	data_out_4,
	data_out_3,
	data_out_2,
	data_out_1,
	data_out_23,
	data_out_22,
	data_out_21,
	data_out_20,
	data_out_19,
	data_out_18,
	data_out_17,
	data_out_16,
	data_out_15,
	data_out_14,
	data_out_13,
	data_valid,
	out_valid,
	out_data_21,
	out_data_20,
	out_data_19,
	out_data_18,
	out_data_17,
	out_data_16,
	out_data_15,
	out_data_14,
	out_data_12,
	out_data_13,
	out_data_9,
	out_data_8,
	out_data_7,
	out_data_6,
	out_data_5,
	out_data_4,
	out_data_3,
	out_data_2,
	out_data_0,
	out_data_1,
	out_data_11,
	out_data_10,
	out_data_23,
	out_data_22,
	clk)/* synthesis synthesis_greybox=0 */;
input 	reset_n;
output 	data_out_12;
output 	data_out_0;
output 	data_out_11;
output 	data_out_10;
output 	data_out_9;
output 	data_out_8;
output 	data_out_7;
output 	data_out_6;
output 	data_out_5;
output 	data_out_4;
output 	data_out_3;
output 	data_out_2;
output 	data_out_1;
output 	data_out_23;
output 	data_out_22;
output 	data_out_21;
output 	data_out_20;
output 	data_out_19;
output 	data_out_18;
output 	data_out_17;
output 	data_out_16;
output 	data_out_15;
output 	data_out_14;
output 	data_out_13;
output 	data_valid;
input 	out_valid;
input 	out_data_21;
input 	out_data_20;
input 	out_data_19;
input 	out_data_18;
input 	out_data_17;
input 	out_data_16;
input 	out_data_15;
input 	out_data_14;
input 	out_data_12;
input 	out_data_13;
input 	out_data_9;
input 	out_data_8;
input 	out_data_7;
input 	out_data_6;
input 	out_data_5;
input 	out_data_4;
input 	out_data_3;
input 	out_data_2;
input 	out_data_0;
input 	out_data_1;
input 	out_data_11;
input 	out_data_10;
input 	out_data_23;
input 	out_data_22;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



lms_dsp_lms_dsp_fir_compiler_ii_0_ast lms_dsp_fir_compiler_ii_0_ast_inst(
	.reset_n(reset_n),
	.data_out_12(data_out_12),
	.data_out_0(data_out_0),
	.data_out_11(data_out_11),
	.data_out_10(data_out_10),
	.data_out_9(data_out_9),
	.data_out_8(data_out_8),
	.data_out_7(data_out_7),
	.data_out_6(data_out_6),
	.data_out_5(data_out_5),
	.data_out_4(data_out_4),
	.data_out_3(data_out_3),
	.data_out_2(data_out_2),
	.data_out_1(data_out_1),
	.data_out_23(data_out_23),
	.data_out_22(data_out_22),
	.data_out_21(data_out_21),
	.data_out_20(data_out_20),
	.data_out_19(data_out_19),
	.data_out_18(data_out_18),
	.data_out_17(data_out_17),
	.data_out_16(data_out_16),
	.data_out_15(data_out_15),
	.data_out_14(data_out_14),
	.data_out_13(data_out_13),
	.data_valid(data_valid),
	.out_valid(out_valid),
	.out_data_21(out_data_21),
	.out_data_20(out_data_20),
	.out_data_19(out_data_19),
	.out_data_18(out_data_18),
	.out_data_17(out_data_17),
	.out_data_16(out_data_16),
	.out_data_15(out_data_15),
	.out_data_14(out_data_14),
	.out_data_12(out_data_12),
	.out_data_13(out_data_13),
	.out_data_9(out_data_9),
	.out_data_8(out_data_8),
	.out_data_7(out_data_7),
	.out_data_6(out_data_6),
	.out_data_5(out_data_5),
	.out_data_4(out_data_4),
	.out_data_3(out_data_3),
	.out_data_2(out_data_2),
	.out_data_0(out_data_0),
	.out_data_1(out_data_1),
	.out_data_11(out_data_11),
	.out_data_10(out_data_10),
	.out_data_23(out_data_23),
	.out_data_22(out_data_22),
	.clk(clk));

endmodule

module lms_dsp_lms_dsp_fir_compiler_ii_0_ast (
	reset_n,
	data_out_12,
	data_out_0,
	data_out_11,
	data_out_10,
	data_out_9,
	data_out_8,
	data_out_7,
	data_out_6,
	data_out_5,
	data_out_4,
	data_out_3,
	data_out_2,
	data_out_1,
	data_out_23,
	data_out_22,
	data_out_21,
	data_out_20,
	data_out_19,
	data_out_18,
	data_out_17,
	data_out_16,
	data_out_15,
	data_out_14,
	data_out_13,
	data_valid,
	out_valid,
	out_data_21,
	out_data_20,
	out_data_19,
	out_data_18,
	out_data_17,
	out_data_16,
	out_data_15,
	out_data_14,
	out_data_12,
	out_data_13,
	out_data_9,
	out_data_8,
	out_data_7,
	out_data_6,
	out_data_5,
	out_data_4,
	out_data_3,
	out_data_2,
	out_data_0,
	out_data_1,
	out_data_11,
	out_data_10,
	out_data_23,
	out_data_22,
	clk)/* synthesis synthesis_greybox=0 */;
input 	reset_n;
output 	data_out_12;
output 	data_out_0;
output 	data_out_11;
output 	data_out_10;
output 	data_out_9;
output 	data_out_8;
output 	data_out_7;
output 	data_out_6;
output 	data_out_5;
output 	data_out_4;
output 	data_out_3;
output 	data_out_2;
output 	data_out_1;
output 	data_out_23;
output 	data_out_22;
output 	data_out_21;
output 	data_out_20;
output 	data_out_19;
output 	data_out_18;
output 	data_out_17;
output 	data_out_16;
output 	data_out_15;
output 	data_out_14;
output 	data_out_13;
output 	data_valid;
input 	out_valid;
input 	out_data_21;
input 	out_data_20;
input 	out_data_19;
input 	out_data_18;
input 	out_data_17;
input 	out_data_16;
input 	out_data_15;
input 	out_data_14;
input 	out_data_12;
input 	out_data_13;
input 	out_data_9;
input 	out_data_8;
input 	out_data_7;
input 	out_data_6;
input 	out_data_5;
input 	out_data_4;
input 	out_data_3;
input 	out_data_2;
input 	out_data_0;
input 	out_data_1;
input 	out_data_11;
input 	out_data_10;
input 	out_data_23;
input 	out_data_22;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[9]~q ;
wire \real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[9]~q ;
wire \real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[20]~q ;
wire \real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[19]~q ;
wire \real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[18]~q ;
wire \real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[17]~q ;
wire \real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[16]~q ;
wire \real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[15]~q ;
wire \real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[14]~q ;
wire \real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[13]~q ;
wire \real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[12]~q ;
wire \real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[11]~q ;
wire \real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[10]~q ;
wire \real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[20]~q ;
wire \real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[19]~q ;
wire \real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[18]~q ;
wire \real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[17]~q ;
wire \real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[16]~q ;
wire \real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[15]~q ;
wire \real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[14]~q ;
wire \real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[13]~q ;
wire \real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[12]~q ;
wire \real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[11]~q ;
wire \real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[10]~q ;
wire \real_passthrough:hpfircore_core|u0_m0_wo0_oseq_gated_reg_q[0]~q ;


lms_dsp_lms_dsp_fir_compiler_ii_0_rtl_core \real_passthrough:hpfircore_core (
	.u1_m0_wo0_mtree_add4_0_o_9(\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[9]~q ),
	.u0_m0_wo0_mtree_add4_0_o_9(\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[9]~q ),
	.u0_m0_wo0_mtree_add4_0_o_20(\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[20]~q ),
	.u0_m0_wo0_mtree_add4_0_o_19(\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[19]~q ),
	.u0_m0_wo0_mtree_add4_0_o_18(\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[18]~q ),
	.u0_m0_wo0_mtree_add4_0_o_17(\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[17]~q ),
	.u0_m0_wo0_mtree_add4_0_o_16(\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[16]~q ),
	.u0_m0_wo0_mtree_add4_0_o_15(\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[15]~q ),
	.u0_m0_wo0_mtree_add4_0_o_14(\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[14]~q ),
	.u0_m0_wo0_mtree_add4_0_o_13(\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[13]~q ),
	.u0_m0_wo0_mtree_add4_0_o_12(\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[12]~q ),
	.u0_m0_wo0_mtree_add4_0_o_11(\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[11]~q ),
	.u0_m0_wo0_mtree_add4_0_o_10(\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[10]~q ),
	.u1_m0_wo0_mtree_add4_0_o_20(\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[20]~q ),
	.u1_m0_wo0_mtree_add4_0_o_19(\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[19]~q ),
	.u1_m0_wo0_mtree_add4_0_o_18(\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[18]~q ),
	.u1_m0_wo0_mtree_add4_0_o_17(\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[17]~q ),
	.u1_m0_wo0_mtree_add4_0_o_16(\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[16]~q ),
	.u1_m0_wo0_mtree_add4_0_o_15(\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[15]~q ),
	.u1_m0_wo0_mtree_add4_0_o_14(\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[14]~q ),
	.u1_m0_wo0_mtree_add4_0_o_13(\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[13]~q ),
	.u1_m0_wo0_mtree_add4_0_o_12(\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[12]~q ),
	.u1_m0_wo0_mtree_add4_0_o_11(\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[11]~q ),
	.u1_m0_wo0_mtree_add4_0_o_10(\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[10]~q ),
	.areset(reset_n),
	.u0_m0_wo0_oseq_gated_reg_q_0(\real_passthrough:hpfircore_core|u0_m0_wo0_oseq_gated_reg_q[0]~q ),
	.xIn_v({out_valid}),
	.xIn_1({out_data_23,out_data_22,out_data_21,out_data_20,out_data_19,out_data_18,out_data_17,out_data_16,out_data_15,out_data_14,out_data_13,out_data_12}),
	.xIn_0({out_data_11,out_data_10,out_data_9,out_data_8,out_data_7,out_data_6,out_data_5,out_data_4,out_data_3,out_data_2,out_data_1,out_data_0}),
	.clk(clk));

lms_dsp_auk_dspip_avalon_streaming_source_hpfir source(
	.data_in({\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[20]~q ,\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[19]~q ,\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[18]~q ,\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[17]~q ,
\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[16]~q ,\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[15]~q ,\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[14]~q ,\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[13]~q ,
\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[12]~q ,\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[11]~q ,\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[10]~q ,\real_passthrough:hpfircore_core|u1_m0_wo0_mtree_add4_0_o[9]~q ,
\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[20]~q ,\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[19]~q ,\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[18]~q ,\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[17]~q ,
\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[16]~q ,\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[15]~q ,\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[14]~q ,\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[13]~q ,
\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[12]~q ,\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[11]~q ,\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[10]~q ,\real_passthrough:hpfircore_core|u0_m0_wo0_mtree_add4_0_o[9]~q }),
	.reset_n(reset_n),
	.data_out_12(data_out_12),
	.data_out_0(data_out_0),
	.data_out_11(data_out_11),
	.data_out_10(data_out_10),
	.data_out_9(data_out_9),
	.data_out_8(data_out_8),
	.data_out_7(data_out_7),
	.data_out_6(data_out_6),
	.data_out_5(data_out_5),
	.data_out_4(data_out_4),
	.data_out_3(data_out_3),
	.data_out_2(data_out_2),
	.data_out_1(data_out_1),
	.data_out_23(data_out_23),
	.data_out_22(data_out_22),
	.data_out_21(data_out_21),
	.data_out_20(data_out_20),
	.data_out_19(data_out_19),
	.data_out_18(data_out_18),
	.data_out_17(data_out_17),
	.data_out_16(data_out_16),
	.data_out_15(data_out_15),
	.data_out_14(data_out_14),
	.data_out_13(data_out_13),
	.data_valid1(data_valid),
	.source_valid_ctrl(\real_passthrough:hpfircore_core|u0_m0_wo0_oseq_gated_reg_q[0]~q ),
	.clk(clk));

endmodule

module lms_dsp_auk_dspip_avalon_streaming_source_hpfir (
	data_in,
	reset_n,
	data_out_12,
	data_out_0,
	data_out_11,
	data_out_10,
	data_out_9,
	data_out_8,
	data_out_7,
	data_out_6,
	data_out_5,
	data_out_4,
	data_out_3,
	data_out_2,
	data_out_1,
	data_out_23,
	data_out_22,
	data_out_21,
	data_out_20,
	data_out_19,
	data_out_18,
	data_out_17,
	data_out_16,
	data_out_15,
	data_out_14,
	data_out_13,
	data_valid1,
	source_valid_ctrl,
	clk)/* synthesis synthesis_greybox=0 */;
input 	[23:0] data_in;
input 	reset_n;
output 	data_out_12;
output 	data_out_0;
output 	data_out_11;
output 	data_out_10;
output 	data_out_9;
output 	data_out_8;
output 	data_out_7;
output 	data_out_6;
output 	data_out_5;
output 	data_out_4;
output 	data_out_3;
output 	data_out_2;
output 	data_out_1;
output 	data_out_23;
output 	data_out_22;
output 	data_out_21;
output 	data_out_20;
output 	data_out_19;
output 	data_out_18;
output 	data_out_17;
output 	data_out_16;
output 	data_out_15;
output 	data_out_14;
output 	data_out_13;
output 	data_valid1;
input 	source_valid_ctrl;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \data_out[12] (
	.clk(clk),
	.d(data_in[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_12),
	.prn(vcc));
defparam \data_out[12] .is_wysiwyg = "true";
defparam \data_out[12] .power_up = "low";

dffeas \data_out[0] (
	.clk(clk),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[11] (
	.clk(clk),
	.d(data_in[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_11),
	.prn(vcc));
defparam \data_out[11] .is_wysiwyg = "true";
defparam \data_out[11] .power_up = "low";

dffeas \data_out[10] (
	.clk(clk),
	.d(data_in[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_10),
	.prn(vcc));
defparam \data_out[10] .is_wysiwyg = "true";
defparam \data_out[10] .power_up = "low";

dffeas \data_out[9] (
	.clk(clk),
	.d(data_in[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_9),
	.prn(vcc));
defparam \data_out[9] .is_wysiwyg = "true";
defparam \data_out[9] .power_up = "low";

dffeas \data_out[8] (
	.clk(clk),
	.d(data_in[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_8),
	.prn(vcc));
defparam \data_out[8] .is_wysiwyg = "true";
defparam \data_out[8] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[23] (
	.clk(clk),
	.d(data_in[23]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_23),
	.prn(vcc));
defparam \data_out[23] .is_wysiwyg = "true";
defparam \data_out[23] .power_up = "low";

dffeas \data_out[22] (
	.clk(clk),
	.d(data_in[22]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_22),
	.prn(vcc));
defparam \data_out[22] .is_wysiwyg = "true";
defparam \data_out[22] .power_up = "low";

dffeas \data_out[21] (
	.clk(clk),
	.d(data_in[21]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_21),
	.prn(vcc));
defparam \data_out[21] .is_wysiwyg = "true";
defparam \data_out[21] .power_up = "low";

dffeas \data_out[20] (
	.clk(clk),
	.d(data_in[20]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_20),
	.prn(vcc));
defparam \data_out[20] .is_wysiwyg = "true";
defparam \data_out[20] .power_up = "low";

dffeas \data_out[19] (
	.clk(clk),
	.d(data_in[19]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_19),
	.prn(vcc));
defparam \data_out[19] .is_wysiwyg = "true";
defparam \data_out[19] .power_up = "low";

dffeas \data_out[18] (
	.clk(clk),
	.d(data_in[18]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_18),
	.prn(vcc));
defparam \data_out[18] .is_wysiwyg = "true";
defparam \data_out[18] .power_up = "low";

dffeas \data_out[17] (
	.clk(clk),
	.d(data_in[17]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_17),
	.prn(vcc));
defparam \data_out[17] .is_wysiwyg = "true";
defparam \data_out[17] .power_up = "low";

dffeas \data_out[16] (
	.clk(clk),
	.d(data_in[16]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_16),
	.prn(vcc));
defparam \data_out[16] .is_wysiwyg = "true";
defparam \data_out[16] .power_up = "low";

dffeas \data_out[15] (
	.clk(clk),
	.d(data_in[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_15),
	.prn(vcc));
defparam \data_out[15] .is_wysiwyg = "true";
defparam \data_out[15] .power_up = "low";

dffeas \data_out[14] (
	.clk(clk),
	.d(data_in[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_14),
	.prn(vcc));
defparam \data_out[14] .is_wysiwyg = "true";
defparam \data_out[14] .power_up = "low";

dffeas \data_out[13] (
	.clk(clk),
	.d(data_in[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_13),
	.prn(vcc));
defparam \data_out[13] .is_wysiwyg = "true";
defparam \data_out[13] .power_up = "low";

dffeas data_valid(
	.clk(clk),
	.d(source_valid_ctrl),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_valid1),
	.prn(vcc));
defparam data_valid.is_wysiwyg = "true";
defparam data_valid.power_up = "low";

endmodule

module lms_dsp_lms_dsp_fir_compiler_ii_0_rtl_core (
	u1_m0_wo0_mtree_add4_0_o_9,
	u0_m0_wo0_mtree_add4_0_o_9,
	u0_m0_wo0_mtree_add4_0_o_20,
	u0_m0_wo0_mtree_add4_0_o_19,
	u0_m0_wo0_mtree_add4_0_o_18,
	u0_m0_wo0_mtree_add4_0_o_17,
	u0_m0_wo0_mtree_add4_0_o_16,
	u0_m0_wo0_mtree_add4_0_o_15,
	u0_m0_wo0_mtree_add4_0_o_14,
	u0_m0_wo0_mtree_add4_0_o_13,
	u0_m0_wo0_mtree_add4_0_o_12,
	u0_m0_wo0_mtree_add4_0_o_11,
	u0_m0_wo0_mtree_add4_0_o_10,
	u1_m0_wo0_mtree_add4_0_o_20,
	u1_m0_wo0_mtree_add4_0_o_19,
	u1_m0_wo0_mtree_add4_0_o_18,
	u1_m0_wo0_mtree_add4_0_o_17,
	u1_m0_wo0_mtree_add4_0_o_16,
	u1_m0_wo0_mtree_add4_0_o_15,
	u1_m0_wo0_mtree_add4_0_o_14,
	u1_m0_wo0_mtree_add4_0_o_13,
	u1_m0_wo0_mtree_add4_0_o_12,
	u1_m0_wo0_mtree_add4_0_o_11,
	u1_m0_wo0_mtree_add4_0_o_10,
	areset,
	u0_m0_wo0_oseq_gated_reg_q_0,
	xIn_v,
	xIn_1,
	xIn_0,
	clk)/* synthesis synthesis_greybox=0 */;
output 	u1_m0_wo0_mtree_add4_0_o_9;
output 	u0_m0_wo0_mtree_add4_0_o_9;
output 	u0_m0_wo0_mtree_add4_0_o_20;
output 	u0_m0_wo0_mtree_add4_0_o_19;
output 	u0_m0_wo0_mtree_add4_0_o_18;
output 	u0_m0_wo0_mtree_add4_0_o_17;
output 	u0_m0_wo0_mtree_add4_0_o_16;
output 	u0_m0_wo0_mtree_add4_0_o_15;
output 	u0_m0_wo0_mtree_add4_0_o_14;
output 	u0_m0_wo0_mtree_add4_0_o_13;
output 	u0_m0_wo0_mtree_add4_0_o_12;
output 	u0_m0_wo0_mtree_add4_0_o_11;
output 	u0_m0_wo0_mtree_add4_0_o_10;
output 	u1_m0_wo0_mtree_add4_0_o_20;
output 	u1_m0_wo0_mtree_add4_0_o_19;
output 	u1_m0_wo0_mtree_add4_0_o_18;
output 	u1_m0_wo0_mtree_add4_0_o_17;
output 	u1_m0_wo0_mtree_add4_0_o_16;
output 	u1_m0_wo0_mtree_add4_0_o_15;
output 	u1_m0_wo0_mtree_add4_0_o_14;
output 	u1_m0_wo0_mtree_add4_0_o_13;
output 	u1_m0_wo0_mtree_add4_0_o_12;
output 	u1_m0_wo0_mtree_add4_0_o_11;
output 	u1_m0_wo0_mtree_add4_0_o_10;
input 	areset;
output 	u0_m0_wo0_oseq_gated_reg_q_0;
input 	[0:0] xIn_v;
input 	[11:0] xIn_1;
input 	[11:0] xIn_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \d_u0_m0_wo0_compute_q_16|delay_signals[0][0]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][9]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][8]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][7]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][6]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][5]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][4]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][3]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][2]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][1]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][0]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][9]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][8]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][7]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][6]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][5]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][4]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][3]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][2]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][1]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][0]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][9]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][8]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][7]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][6]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][5]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][4]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][3]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][2]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][1]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][0]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][9]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][8]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][7]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][6]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][5]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][4]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][3]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][2]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][1]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][0]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][11]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][10]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][11]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][10]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][11]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][10]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][11]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][0]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][9]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][8]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][7]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][6]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][5]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][4]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][3]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][2]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][0]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][0]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][9]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][8]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][7]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][6]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][5]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][4]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][3]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][2]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][0]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][10]~q ;
wire \u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][10]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][11]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][10]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][11]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][10]~q ;
wire \d_u0_m0_wo0_compute_q_13|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][0]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][7]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][6]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][5]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][4]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][3]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][2]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][1]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][6]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][5]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][4]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][3]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][2]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][1]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][7]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][9]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][6]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][8]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][5]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][4]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][3]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][2]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][1]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][0]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][7]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][6]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][5]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][4]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][3]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][2]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][1]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][6]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][5]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][4]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][3]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][2]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][1]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][7]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][9]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][6]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][8]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][5]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][4]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][3]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][2]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][1]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][10]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][11]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][10]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][9]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][8]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][11]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][10]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][9]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][8]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][7]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][10]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][10]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][11]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][10]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][9]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][8]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][11]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][10]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][9]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][8]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][7]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][10]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][11]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][9]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][8]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][7]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][6]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][5]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][4]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][3]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][2]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][1]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][6]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][5]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][4]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][3]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][2]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][1]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][4]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][3]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][2]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][1]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][4]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][3]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][2]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][2]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][9]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][1]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][8]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][0]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][7]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][6]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][5]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][4]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][3]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][4]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][3]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][2]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][4]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][3]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][2]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][1]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][6]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][8]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][9]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][7]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][5]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][4]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][3]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][2]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][1]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][0]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][7]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][6]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][5]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][4]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][3]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][2]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][1]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][8]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][7]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][6]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][5]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][4]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][3]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][2]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][1]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][0]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][9]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][8]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][7]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][6]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][5]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][4]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][3]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][2]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][1]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][6]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][5]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][4]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][3]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][2]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][1]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][4]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][3]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][2]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][1]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][4]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][3]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][2]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][2]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][9]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][1]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][8]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][0]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][7]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][6]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][5]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][4]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][3]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][4]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][3]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][2]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][4]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][3]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][2]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][1]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][6]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][8]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][9]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][7]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][5]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][4]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][3]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][2]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][1]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][0]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][7]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][6]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][5]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][4]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][3]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][2]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][1]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][8]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][7]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][6]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][5]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][4]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][3]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][2]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][1]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][0]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][11]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][10]~q ;
wire \u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][10]~q ;
wire \u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][10]~q ;
wire \u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][10]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][11]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][10]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][9]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][8]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][7]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][11]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][10]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][9]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][8]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][7]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][6]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][5]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][11]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][10]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][9]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][8]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][7]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][6]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][5]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][10]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][11]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][11]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][10]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][9]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][8]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][7]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][6]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][5]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][11]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][10]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][9]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][8]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][7]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][6]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][5]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][11]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][10]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][11]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][10]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][9]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][8]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][11]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][10]~q ;
wire \d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][9]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][11]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][10]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][11]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][10]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][9]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][8]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][7]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][11]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][10]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][9]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][8]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][7]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][6]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][5]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][11]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][10]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][9]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][8]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][7]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][6]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][5]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][10]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][11]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][11]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][10]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][9]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][8]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][7]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][6]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][5]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][11]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][10]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][9]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][8]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][7]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][6]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][5]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][11]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][10]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][11]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][10]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][9]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][8]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][11]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][10]~q ;
wire \d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][9]~q ;
wire \d_u0_m0_wo0_compute_q_11|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][10]~q ;
wire \u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][10]~q ;
wire \u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][10]~q ;
wire \u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][10]~q ;
wire \u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][10]~q ;
wire \u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][10]~q ;
wire \u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][10]~q ;
wire \u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][10]~q ;
wire \u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][10]~q ;
wire \u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][10]~q ;
wire \u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][10]~q ;
wire \u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][10]~q ;
wire \u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][1]~q ;
wire \u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][10]~q ;
wire \u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][10]~q ;
wire \u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][9]~q ;
wire \u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][8]~q ;
wire \u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][7]~q ;
wire \u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][6]~q ;
wire \u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][5]~q ;
wire \u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][4]~q ;
wire \u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][3]~q ;
wire \u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][2]~q ;
wire \u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][0]~q ;
wire \u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][9]~q ;
wire \u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][8]~q ;
wire \u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][7]~q ;
wire \u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][6]~q ;
wire \u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][5]~q ;
wire \u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][4]~q ;
wire \u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][3]~q ;
wire \u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][2]~q ;
wire \u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][0]~q ;
wire \u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][1]~q ;
wire \u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][11]~q ;
wire \u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][10]~q ;
wire \u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][11]~q ;
wire \u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][10]~q ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[1]~13 ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[2]~15 ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[3]~17 ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[4]~19 ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[5]~21 ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[6]~23 ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[7]~25 ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[8]~27 ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[9]~28_combout ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[8]~26_combout ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[7]~24_combout ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[6]~22_combout ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[5]~20_combout ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[4]~18_combout ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[3]~16_combout ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[2]~14_combout ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[1]~12_combout ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[0]~q ;
wire \u1_m0_wo0_mtree_add1_1_o[0]~15 ;
wire \u1_m0_wo0_mtree_add1_1_o[1]~17 ;
wire \u1_m0_wo0_mtree_add1_1_o[2]~19 ;
wire \u1_m0_wo0_mtree_add1_1_o[3]~21 ;
wire \u1_m0_wo0_mtree_add1_1_o[4]~23 ;
wire \u1_m0_wo0_mtree_add1_1_o[5]~25 ;
wire \u1_m0_wo0_mtree_add1_1_o[6]~27 ;
wire \u1_m0_wo0_mtree_add1_1_o[7]~29 ;
wire \u1_m0_wo0_mtree_add1_1_o[8]~31 ;
wire \u1_m0_wo0_mtree_add1_1_o[9]~32_combout ;
wire \u1_m0_wo0_mtree_add1_1_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[2]~14 ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[3]~16 ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[4]~18 ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[5]~20 ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[6]~22 ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[7]~24 ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[8]~26 ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[9]~27_combout ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[1]~14 ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[2]~16 ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[3]~18 ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[4]~20 ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[5]~22 ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[6]~24 ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[7]~26 ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[8]~27_combout ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[8]~25_combout ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[7]~25_combout ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[7]~23_combout ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[6]~23_combout ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[6]~21_combout ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[5]~21_combout ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[5]~19_combout ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[4]~19_combout ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[4]~17_combout ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[3]~17_combout ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[3]~15_combout ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[2]~15_combout ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[2]~13_combout ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[1]~13_combout ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[0]~q ;
wire \u1_m0_wo0_mtree_add0_4_o[1]~16 ;
wire \u1_m0_wo0_mtree_add0_4_o[2]~18 ;
wire \u1_m0_wo0_mtree_add0_4_o[3]~20 ;
wire \u1_m0_wo0_mtree_add0_4_o[4]~22 ;
wire \u1_m0_wo0_mtree_add0_4_o[5]~24 ;
wire \u1_m0_wo0_mtree_add0_4_o[6]~26 ;
wire \u1_m0_wo0_mtree_add0_4_o[7]~28 ;
wire \u1_m0_wo0_mtree_add0_4_o[8]~30 ;
wire \u1_m0_wo0_mtree_add0_4_o[9]~31_combout ;
wire \u1_m0_wo0_mtree_add0_4_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[1]~13 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[2]~15 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[3]~17 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[4]~19 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[5]~21 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[6]~23 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[7]~25 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[8]~27 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[9]~28_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[8]~26_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[7]~24_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[6]~22_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[5]~20_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[4]~18_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[3]~16_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[0]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[2]~14_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[2]~14 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[3]~16 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[4]~18 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[5]~20 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[6]~22 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[7]~24 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[8]~26 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[9]~27_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[9]~q ;
wire \u1_m0_wo0_mtree_add0_4_o[8]~29_combout ;
wire \u1_m0_wo0_mtree_add0_4_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[8]~25_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[8]~q ;
wire \u1_m0_wo0_mtree_add0_4_o[7]~27_combout ;
wire \u1_m0_wo0_mtree_add0_4_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[7]~23_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[7]~q ;
wire \u1_m0_wo0_mtree_add0_4_o[6]~25_combout ;
wire \u1_m0_wo0_mtree_add0_4_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[6]~21_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[6]~q ;
wire \u1_m0_wo0_mtree_add0_4_o[5]~23_combout ;
wire \u1_m0_wo0_mtree_add0_4_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[5]~19_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[5]~q ;
wire \u1_m0_wo0_mtree_add0_4_o[4]~21_combout ;
wire \u1_m0_wo0_mtree_add0_4_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[4]~17_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[4]~q ;
wire \u1_m0_wo0_mtree_add0_4_o[3]~19_combout ;
wire \u1_m0_wo0_mtree_add0_4_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[3]~15_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[3]~q ;
wire \u1_m0_wo0_mtree_add0_4_o[2]~17_combout ;
wire \u1_m0_wo0_mtree_add0_4_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[2]~13_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[2]~q ;
wire \u1_m0_wo0_mtree_add0_4_o[1]~15_combout ;
wire \u1_m0_wo0_mtree_add0_4_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[1]~12_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[0]~q ;
wire \u1_m0_wo0_mtree_add0_4_o[0]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[0]~q ;
wire \u1_m0_wo0_mtree_add1_2_o[0]~18 ;
wire \u1_m0_wo0_mtree_add1_2_o[1]~20 ;
wire \u1_m0_wo0_mtree_add1_2_o[2]~22 ;
wire \u1_m0_wo0_mtree_add1_2_o[3]~24 ;
wire \u1_m0_wo0_mtree_add1_2_o[4]~26 ;
wire \u1_m0_wo0_mtree_add1_2_o[5]~28 ;
wire \u1_m0_wo0_mtree_add1_2_o[6]~30 ;
wire \u1_m0_wo0_mtree_add1_2_o[7]~32 ;
wire \u1_m0_wo0_mtree_add1_2_o[8]~34 ;
wire \u1_m0_wo0_mtree_add1_2_o[9]~35_combout ;
wire \u1_m0_wo0_mtree_add1_2_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[1]~14 ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[2]~16 ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[3]~18 ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[4]~20 ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[5]~22 ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[6]~24 ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[7]~26 ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[8]~28 ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[9]~29_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[8]~27_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[7]~25_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[6]~23_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[5]~21_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[4]~19_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[0]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[3]~17_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[3]~14 ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[4]~16 ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[5]~18 ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[6]~20 ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[7]~22 ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[8]~24 ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[9]~25_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[1]~16 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[2]~18 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[3]~20 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[4]~22 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[5]~24 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[6]~26 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[7]~28 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[8]~30 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[9]~31_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[8]~29_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[7]~27_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[6]~25_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[0]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[5]~23_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[5]~14 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[6]~16 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[7]~18 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[8]~20 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[9]~21_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[8]~23_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[8]~19_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[7]~21_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[7]~17_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[6]~19_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[6]~15_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[5]~17_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[5]~13_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[4]~15_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[4]~21_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[3]~13_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[3]~19_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[2]~15_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[2]~17_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[1]~13_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[1]~15_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[0]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[0]~q ;
wire \u1_m0_wo0_mtree_add0_6_o[0]~20 ;
wire \u1_m0_wo0_mtree_add0_6_o[1]~22 ;
wire \u1_m0_wo0_mtree_add0_6_o[2]~24 ;
wire \u1_m0_wo0_mtree_add0_6_o[3]~26 ;
wire \u1_m0_wo0_mtree_add0_6_o[4]~28 ;
wire \u1_m0_wo0_mtree_add0_6_o[5]~30 ;
wire \u1_m0_wo0_mtree_add0_6_o[6]~32 ;
wire \u1_m0_wo0_mtree_add0_6_o[7]~34 ;
wire \u1_m0_wo0_mtree_add0_6_o[8]~36 ;
wire \u1_m0_wo0_mtree_add0_6_o[9]~37_combout ;
wire \u1_m0_wo0_mtree_add0_6_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[2]~14 ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[3]~16 ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[4]~18 ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[5]~20 ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[6]~22 ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[7]~24 ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[8]~26 ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[9]~27_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[8]~25_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[7]~23_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[6]~21_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[0]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[5]~19_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[5]~14 ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[6]~16 ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[7]~18 ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[8]~20 ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[9]~21_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[1]~20 ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[2]~22 ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[3]~24 ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[4]~26 ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[5]~28 ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[6]~30 ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[7]~32 ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[8]~34 ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[9]~35_combout ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[8]~19_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[8]~33_combout ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[7]~17_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[7]~31_combout ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[6]~15_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[6]~29_combout ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[5]~13_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[5]~27_combout ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[4]~17_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[4]~25_combout ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[3]~15_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[3]~23_combout ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[2]~13_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[2]~21_combout ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[1]~19_combout ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[0]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[0]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[0]~22 ;
wire \u1_m0_wo0_mtree_add0_7_o[1]~24 ;
wire \u1_m0_wo0_mtree_add0_7_o[2]~26 ;
wire \u1_m0_wo0_mtree_add0_7_o[3]~28 ;
wire \u1_m0_wo0_mtree_add0_7_o[4]~30 ;
wire \u1_m0_wo0_mtree_add0_7_o[5]~32 ;
wire \u1_m0_wo0_mtree_add0_7_o[6]~34 ;
wire \u1_m0_wo0_mtree_add0_7_o[7]~36 ;
wire \u1_m0_wo0_mtree_add0_7_o[8]~38 ;
wire \u1_m0_wo0_mtree_add0_7_o[9]~39_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[9]~q ;
wire \u1_m0_wo0_mtree_add0_6_o[8]~35_combout ;
wire \u1_m0_wo0_mtree_add0_6_o[8]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[8]~37_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[8]~q ;
wire \u1_m0_wo0_mtree_add0_6_o[7]~33_combout ;
wire \u1_m0_wo0_mtree_add0_6_o[7]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[7]~35_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[7]~q ;
wire \u1_m0_wo0_mtree_add0_6_o[6]~31_combout ;
wire \u1_m0_wo0_mtree_add0_6_o[6]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[6]~33_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[6]~q ;
wire \u1_m0_wo0_mtree_add0_6_o[5]~29_combout ;
wire \u1_m0_wo0_mtree_add0_6_o[5]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[5]~31_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[5]~q ;
wire \u1_m0_wo0_mtree_add0_6_o[4]~27_combout ;
wire \u1_m0_wo0_mtree_add0_6_o[4]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[4]~29_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[4]~q ;
wire \u1_m0_wo0_mtree_add0_6_o[3]~25_combout ;
wire \u1_m0_wo0_mtree_add0_6_o[3]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[3]~27_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[3]~q ;
wire \u1_m0_wo0_mtree_add0_6_o[2]~23_combout ;
wire \u1_m0_wo0_mtree_add0_6_o[2]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[2]~25_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[2]~q ;
wire \u1_m0_wo0_mtree_add0_6_o[1]~21_combout ;
wire \u1_m0_wo0_mtree_add0_6_o[1]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[1]~23_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[1]~q ;
wire \u1_m0_wo0_mtree_add0_6_o[0]~19_combout ;
wire \u1_m0_wo0_mtree_add0_6_o[0]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[0]~21_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[0]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[0]~22 ;
wire \u1_m0_wo0_mtree_add1_3_o[1]~24 ;
wire \u1_m0_wo0_mtree_add1_3_o[2]~26 ;
wire \u1_m0_wo0_mtree_add1_3_o[3]~28 ;
wire \u1_m0_wo0_mtree_add1_3_o[4]~30 ;
wire \u1_m0_wo0_mtree_add1_3_o[5]~32 ;
wire \u1_m0_wo0_mtree_add1_3_o[6]~34 ;
wire \u1_m0_wo0_mtree_add1_3_o[7]~36 ;
wire \u1_m0_wo0_mtree_add1_3_o[8]~38 ;
wire \u1_m0_wo0_mtree_add1_3_o[9]~39_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[9]~q ;
wire \u1_m0_wo0_mtree_add1_2_o[8]~33_combout ;
wire \u1_m0_wo0_mtree_add1_2_o[8]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[8]~37_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[8]~q ;
wire \u1_m0_wo0_mtree_add1_2_o[7]~31_combout ;
wire \u1_m0_wo0_mtree_add1_2_o[7]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[7]~35_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[7]~q ;
wire \u1_m0_wo0_mtree_add1_2_o[6]~29_combout ;
wire \u1_m0_wo0_mtree_add1_2_o[6]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[6]~33_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[6]~q ;
wire \u1_m0_wo0_mtree_add1_2_o[5]~27_combout ;
wire \u1_m0_wo0_mtree_add1_2_o[5]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[5]~31_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[5]~q ;
wire \u1_m0_wo0_mtree_add1_2_o[4]~25_combout ;
wire \u1_m0_wo0_mtree_add1_2_o[4]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[4]~29_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[4]~q ;
wire \u1_m0_wo0_mtree_add1_2_o[3]~23_combout ;
wire \u1_m0_wo0_mtree_add1_2_o[3]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[3]~27_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[3]~q ;
wire \u1_m0_wo0_mtree_add1_2_o[2]~21_combout ;
wire \u1_m0_wo0_mtree_add1_2_o[2]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[2]~25_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[2]~q ;
wire \u1_m0_wo0_mtree_add1_2_o[1]~19_combout ;
wire \u1_m0_wo0_mtree_add1_2_o[1]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[1]~23_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[1]~q ;
wire \u1_m0_wo0_mtree_add1_2_o[0]~17_combout ;
wire \u1_m0_wo0_mtree_add1_2_o[0]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[0]~21_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[0]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[0]~22 ;
wire \u1_m0_wo0_mtree_add2_1_o[1]~24 ;
wire \u1_m0_wo0_mtree_add2_1_o[2]~26 ;
wire \u1_m0_wo0_mtree_add2_1_o[3]~28 ;
wire \u1_m0_wo0_mtree_add2_1_o[4]~30 ;
wire \u1_m0_wo0_mtree_add2_1_o[5]~32 ;
wire \u1_m0_wo0_mtree_add2_1_o[6]~34 ;
wire \u1_m0_wo0_mtree_add2_1_o[7]~36 ;
wire \u1_m0_wo0_mtree_add2_1_o[8]~38 ;
wire \u1_m0_wo0_mtree_add2_1_o[9]~39_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[9]~q ;
wire \u1_m0_wo0_mtree_add1_1_o[8]~30_combout ;
wire \u1_m0_wo0_mtree_add1_1_o[8]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[8]~37_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[8]~q ;
wire \u1_m0_wo0_mtree_add1_1_o[7]~28_combout ;
wire \u1_m0_wo0_mtree_add1_1_o[7]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[7]~35_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[7]~q ;
wire \u1_m0_wo0_mtree_add1_1_o[6]~26_combout ;
wire \u1_m0_wo0_mtree_add1_1_o[6]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[6]~33_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[6]~q ;
wire \u1_m0_wo0_mtree_add1_1_o[5]~24_combout ;
wire \u1_m0_wo0_mtree_add1_1_o[5]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[5]~31_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[5]~q ;
wire \u1_m0_wo0_mtree_add1_1_o[4]~22_combout ;
wire \u1_m0_wo0_mtree_add1_1_o[4]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[4]~29_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[4]~q ;
wire \u1_m0_wo0_mtree_add1_1_o[3]~20_combout ;
wire \u1_m0_wo0_mtree_add1_1_o[3]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[3]~27_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[3]~q ;
wire \u1_m0_wo0_mtree_add1_1_o[2]~18_combout ;
wire \u1_m0_wo0_mtree_add1_1_o[2]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[2]~25_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[2]~q ;
wire \u1_m0_wo0_mtree_add1_1_o[1]~16_combout ;
wire \u1_m0_wo0_mtree_add1_1_o[1]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[1]~23_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[1]~q ;
wire \u1_m0_wo0_mtree_add1_1_o[0]~14_combout ;
wire \u1_m0_wo0_mtree_add1_1_o[0]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[0]~21_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[0]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[0]~22 ;
wire \u1_m0_wo0_mtree_add3_0_o[1]~24 ;
wire \u1_m0_wo0_mtree_add3_0_o[2]~26 ;
wire \u1_m0_wo0_mtree_add3_0_o[3]~28 ;
wire \u1_m0_wo0_mtree_add3_0_o[4]~30 ;
wire \u1_m0_wo0_mtree_add3_0_o[5]~32 ;
wire \u1_m0_wo0_mtree_add3_0_o[6]~34 ;
wire \u1_m0_wo0_mtree_add3_0_o[7]~36 ;
wire \u1_m0_wo0_mtree_add3_0_o[8]~38 ;
wire \u1_m0_wo0_mtree_add3_0_o[9]~39_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[2]~14 ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[3]~16 ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[4]~18 ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[5]~20 ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[6]~22 ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[7]~24 ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[8]~26 ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[9]~27_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[8]~25_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[7]~23_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[6]~21_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[0]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[5]~19_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[5]~14 ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[6]~16 ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[7]~18 ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[8]~20 ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[9]~21_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[1]~16 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[2]~18 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[3]~20 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[4]~22 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[5]~24 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[6]~26 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[7]~28 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[8]~30 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[9]~31_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[8]~29_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[7]~27_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[6]~25_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[0]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[5]~23_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[5]~14 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[6]~16 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[7]~18 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[8]~20 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[9]~21_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[8]~19_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[8]~19_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[7]~17_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[7]~17_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[6]~15_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[6]~15_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[5]~13_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[5]~13_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[4]~17_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[4]~21_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[3]~15_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[3]~19_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[2]~13_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[2]~17_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[1]~15_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[0]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[0]~q ;
wire \u1_m0_wo0_mtree_add0_8_o[0]~20 ;
wire \u1_m0_wo0_mtree_add0_8_o[1]~22 ;
wire \u1_m0_wo0_mtree_add0_8_o[2]~24 ;
wire \u1_m0_wo0_mtree_add0_8_o[3]~26 ;
wire \u1_m0_wo0_mtree_add0_8_o[4]~28 ;
wire \u1_m0_wo0_mtree_add0_8_o[5]~30 ;
wire \u1_m0_wo0_mtree_add0_8_o[6]~32 ;
wire \u1_m0_wo0_mtree_add0_8_o[7]~34 ;
wire \u1_m0_wo0_mtree_add0_8_o[8]~36 ;
wire \u1_m0_wo0_mtree_add0_8_o[9]~37_combout ;
wire \u1_m0_wo0_mtree_add0_8_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[1]~14 ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[2]~16 ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[3]~18 ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[4]~20 ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[5]~22 ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[6]~24 ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[7]~26 ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[8]~28 ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[9]~29_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[8]~27_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[7]~25_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[6]~23_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[5]~21_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[4]~19_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[0]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[3]~17_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[3]~14 ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[4]~16 ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[5]~18 ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[6]~20 ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[7]~22 ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[8]~24 ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[9]~25_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[9]~q ;
wire \u1_m0_wo0_mtree_add0_8_o[8]~35_combout ;
wire \u1_m0_wo0_mtree_add0_8_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[8]~23_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[8]~q ;
wire \u1_m0_wo0_mtree_add0_8_o[7]~33_combout ;
wire \u1_m0_wo0_mtree_add0_8_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[7]~21_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[7]~q ;
wire \u1_m0_wo0_mtree_add0_8_o[6]~31_combout ;
wire \u1_m0_wo0_mtree_add0_8_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[6]~19_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[6]~q ;
wire \u1_m0_wo0_mtree_add0_8_o[5]~29_combout ;
wire \u1_m0_wo0_mtree_add0_8_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[5]~17_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[5]~q ;
wire \u1_m0_wo0_mtree_add0_8_o[4]~27_combout ;
wire \u1_m0_wo0_mtree_add0_8_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[4]~15_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[4]~q ;
wire \u1_m0_wo0_mtree_add0_8_o[3]~25_combout ;
wire \u1_m0_wo0_mtree_add0_8_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[3]~13_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[3]~q ;
wire \u1_m0_wo0_mtree_add0_8_o[2]~23_combout ;
wire \u1_m0_wo0_mtree_add0_8_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[2]~15_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[2]~q ;
wire \u1_m0_wo0_mtree_add0_8_o[1]~21_combout ;
wire \u1_m0_wo0_mtree_add0_8_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[1]~13_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[1]~q ;
wire \u1_m0_wo0_mtree_add0_8_o[0]~19_combout ;
wire \u1_m0_wo0_mtree_add0_8_o[0]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[0]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[0]~21 ;
wire \u1_m0_wo0_mtree_add1_4_o[1]~23 ;
wire \u1_m0_wo0_mtree_add1_4_o[2]~25 ;
wire \u1_m0_wo0_mtree_add1_4_o[3]~27 ;
wire \u1_m0_wo0_mtree_add1_4_o[4]~29 ;
wire \u1_m0_wo0_mtree_add1_4_o[5]~31 ;
wire \u1_m0_wo0_mtree_add1_4_o[6]~33 ;
wire \u1_m0_wo0_mtree_add1_4_o[7]~35 ;
wire \u1_m0_wo0_mtree_add1_4_o[8]~37 ;
wire \u1_m0_wo0_mtree_add1_4_o[9]~38_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[1]~13 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[2]~15 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[3]~17 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[4]~19 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[5]~21 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[6]~23 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[7]~25 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[8]~27 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[9]~28_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[8]~26_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[7]~24_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[6]~22_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[5]~20_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[4]~18_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[3]~16_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[0]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[2]~14_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[2]~14 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[3]~16 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[4]~18 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[5]~20 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[6]~22 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[7]~24 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[8]~26 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[9]~27_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[1]~14 ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[2]~16 ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[3]~18 ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[4]~20 ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[5]~22 ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[6]~24 ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[7]~26 ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[8]~27_combout ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[8]~25_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[7]~25_combout ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[7]~23_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[6]~23_combout ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[6]~21_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[5]~21_combout ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[5]~19_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[4]~19_combout ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[4]~17_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[3]~17_combout ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[3]~15_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[2]~15_combout ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[2]~13_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[1]~13_combout ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[1]~12_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[0]~q ;
wire \u1_m0_wo0_mtree_add0_10_o[1]~16 ;
wire \u1_m0_wo0_mtree_add0_10_o[2]~18 ;
wire \u1_m0_wo0_mtree_add0_10_o[3]~20 ;
wire \u1_m0_wo0_mtree_add0_10_o[4]~22 ;
wire \u1_m0_wo0_mtree_add0_10_o[5]~24 ;
wire \u1_m0_wo0_mtree_add0_10_o[6]~26 ;
wire \u1_m0_wo0_mtree_add0_10_o[7]~28 ;
wire \u1_m0_wo0_mtree_add0_10_o[8]~30 ;
wire \u1_m0_wo0_mtree_add0_10_o[9]~31_combout ;
wire \u1_m0_wo0_mtree_add0_10_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[2]~14 ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[3]~16 ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[4]~18 ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[5]~20 ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[6]~22 ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[7]~24 ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[8]~26 ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[9]~27_combout ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[9]~q ;
wire \u1_m0_wo0_mtree_add0_10_o[8]~29_combout ;
wire \u1_m0_wo0_mtree_add0_10_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[8]~25_combout ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[8]~q ;
wire \u1_m0_wo0_mtree_add0_10_o[7]~27_combout ;
wire \u1_m0_wo0_mtree_add0_10_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[7]~23_combout ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[7]~q ;
wire \u1_m0_wo0_mtree_add0_10_o[6]~25_combout ;
wire \u1_m0_wo0_mtree_add0_10_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[6]~21_combout ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[6]~q ;
wire \u1_m0_wo0_mtree_add0_10_o[5]~23_combout ;
wire \u1_m0_wo0_mtree_add0_10_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[5]~19_combout ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[5]~q ;
wire \u1_m0_wo0_mtree_add0_10_o[4]~21_combout ;
wire \u1_m0_wo0_mtree_add0_10_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[4]~17_combout ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[4]~q ;
wire \u1_m0_wo0_mtree_add0_10_o[3]~19_combout ;
wire \u1_m0_wo0_mtree_add0_10_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[3]~15_combout ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[3]~q ;
wire \u1_m0_wo0_mtree_add0_10_o[2]~17_combout ;
wire \u1_m0_wo0_mtree_add0_10_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[2]~13_combout ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[2]~q ;
wire \u1_m0_wo0_mtree_add0_10_o[1]~15_combout ;
wire \u1_m0_wo0_mtree_add0_10_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[0]~q ;
wire \u1_m0_wo0_mtree_add0_10_o[0]~q ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[0]~q ;
wire \u1_m0_wo0_mtree_add1_5_o[0]~18 ;
wire \u1_m0_wo0_mtree_add1_5_o[1]~20 ;
wire \u1_m0_wo0_mtree_add1_5_o[2]~22 ;
wire \u1_m0_wo0_mtree_add1_5_o[3]~24 ;
wire \u1_m0_wo0_mtree_add1_5_o[4]~26 ;
wire \u1_m0_wo0_mtree_add1_5_o[5]~28 ;
wire \u1_m0_wo0_mtree_add1_5_o[6]~30 ;
wire \u1_m0_wo0_mtree_add1_5_o[7]~32 ;
wire \u1_m0_wo0_mtree_add1_5_o[8]~34 ;
wire \u1_m0_wo0_mtree_add1_5_o[9]~35_combout ;
wire \u1_m0_wo0_mtree_add1_5_o[9]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[8]~36_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[8]~q ;
wire \u1_m0_wo0_mtree_add1_5_o[8]~33_combout ;
wire \u1_m0_wo0_mtree_add1_5_o[8]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[7]~34_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[7]~q ;
wire \u1_m0_wo0_mtree_add1_5_o[7]~31_combout ;
wire \u1_m0_wo0_mtree_add1_5_o[7]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[6]~32_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[6]~q ;
wire \u1_m0_wo0_mtree_add1_5_o[6]~29_combout ;
wire \u1_m0_wo0_mtree_add1_5_o[6]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[5]~30_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[5]~q ;
wire \u1_m0_wo0_mtree_add1_5_o[5]~27_combout ;
wire \u1_m0_wo0_mtree_add1_5_o[5]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[4]~28_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[4]~q ;
wire \u1_m0_wo0_mtree_add1_5_o[4]~25_combout ;
wire \u1_m0_wo0_mtree_add1_5_o[4]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[3]~26_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[3]~q ;
wire \u1_m0_wo0_mtree_add1_5_o[3]~23_combout ;
wire \u1_m0_wo0_mtree_add1_5_o[3]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[2]~24_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[2]~q ;
wire \u1_m0_wo0_mtree_add1_5_o[2]~21_combout ;
wire \u1_m0_wo0_mtree_add1_5_o[2]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[1]~22_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[1]~q ;
wire \u1_m0_wo0_mtree_add1_5_o[1]~19_combout ;
wire \u1_m0_wo0_mtree_add1_5_o[1]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[0]~20_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[0]~q ;
wire \u1_m0_wo0_mtree_add1_5_o[0]~17_combout ;
wire \u1_m0_wo0_mtree_add1_5_o[0]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[0]~22 ;
wire \u1_m0_wo0_mtree_add2_2_o[1]~24 ;
wire \u1_m0_wo0_mtree_add2_2_o[2]~26 ;
wire \u1_m0_wo0_mtree_add2_2_o[3]~28 ;
wire \u1_m0_wo0_mtree_add2_2_o[4]~30 ;
wire \u1_m0_wo0_mtree_add2_2_o[5]~32 ;
wire \u1_m0_wo0_mtree_add2_2_o[6]~34 ;
wire \u1_m0_wo0_mtree_add2_2_o[7]~36 ;
wire \u1_m0_wo0_mtree_add2_2_o[8]~38 ;
wire \u1_m0_wo0_mtree_add2_2_o[9]~39_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[1]~13 ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[2]~15 ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[3]~17 ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[4]~19 ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[5]~21 ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[6]~23 ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[7]~25 ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[8]~27 ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[9]~28_combout ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[9]~q ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[8]~26_combout ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[8]~q ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[7]~24_combout ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[7]~q ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[6]~22_combout ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[6]~q ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[5]~20_combout ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[5]~q ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[4]~18_combout ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[4]~q ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[3]~16_combout ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[3]~q ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[2]~14_combout ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[2]~q ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[1]~12_combout ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[1]~q ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[0]~q ;
wire \u1_m0_wo0_mtree_add0_12_o[0]~15 ;
wire \u1_m0_wo0_mtree_add0_12_o[1]~17 ;
wire \u1_m0_wo0_mtree_add0_12_o[2]~19 ;
wire \u1_m0_wo0_mtree_add0_12_o[3]~21 ;
wire \u1_m0_wo0_mtree_add0_12_o[4]~23 ;
wire \u1_m0_wo0_mtree_add0_12_o[5]~25 ;
wire \u1_m0_wo0_mtree_add0_12_o[6]~27 ;
wire \u1_m0_wo0_mtree_add0_12_o[7]~29 ;
wire \u1_m0_wo0_mtree_add0_12_o[8]~31 ;
wire \u1_m0_wo0_mtree_add0_12_o[9]~32_combout ;
wire \u1_m0_wo0_mtree_add0_12_o[9]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[8]~37_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[8]~q ;
wire \u1_m0_wo0_mtree_add0_12_o[8]~30_combout ;
wire \u1_m0_wo0_mtree_add0_12_o[8]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[7]~35_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[7]~q ;
wire \u1_m0_wo0_mtree_add0_12_o[7]~28_combout ;
wire \u1_m0_wo0_mtree_add0_12_o[7]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[6]~33_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[6]~q ;
wire \u1_m0_wo0_mtree_add0_12_o[6]~26_combout ;
wire \u1_m0_wo0_mtree_add0_12_o[6]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[5]~31_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[5]~q ;
wire \u1_m0_wo0_mtree_add0_12_o[5]~24_combout ;
wire \u1_m0_wo0_mtree_add0_12_o[5]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[4]~29_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[4]~q ;
wire \u1_m0_wo0_mtree_add0_12_o[4]~22_combout ;
wire \u1_m0_wo0_mtree_add0_12_o[4]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[3]~27_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[3]~q ;
wire \u1_m0_wo0_mtree_add0_12_o[3]~20_combout ;
wire \u1_m0_wo0_mtree_add0_12_o[3]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[2]~25_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[2]~q ;
wire \u1_m0_wo0_mtree_add0_12_o[2]~18_combout ;
wire \u1_m0_wo0_mtree_add0_12_o[2]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[1]~23_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[1]~q ;
wire \u1_m0_wo0_mtree_add0_12_o[1]~16_combout ;
wire \u1_m0_wo0_mtree_add0_12_o[1]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[0]~21_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[0]~q ;
wire \u1_m0_wo0_mtree_add0_12_o[0]~14_combout ;
wire \u1_m0_wo0_mtree_add0_12_o[0]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[0]~22 ;
wire \u1_m0_wo0_mtree_add3_1_o[1]~24 ;
wire \u1_m0_wo0_mtree_add3_1_o[2]~26 ;
wire \u1_m0_wo0_mtree_add3_1_o[3]~28 ;
wire \u1_m0_wo0_mtree_add3_1_o[4]~30 ;
wire \u1_m0_wo0_mtree_add3_1_o[5]~32 ;
wire \u1_m0_wo0_mtree_add3_1_o[6]~34 ;
wire \u1_m0_wo0_mtree_add3_1_o[7]~36 ;
wire \u1_m0_wo0_mtree_add3_1_o[8]~38 ;
wire \u1_m0_wo0_mtree_add3_1_o[9]~39_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[9]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[8]~37_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[8]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[8]~37_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[8]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[7]~35_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[7]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[7]~35_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[7]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[6]~33_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[6]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[6]~33_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[6]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[5]~31_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[5]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[5]~31_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[5]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[4]~29_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[4]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[4]~29_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[4]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[3]~27_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[3]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[3]~27_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[3]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[2]~25_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[2]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[2]~25_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[2]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[1]~23_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[1]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[1]~23_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[1]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[0]~21_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[0]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[0]~21_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[0]~q ;
wire \u1_m0_wo0_mtree_add4_0_o[9]~13_cout ;
wire \u1_m0_wo0_mtree_add4_0_o[9]~15_cout ;
wire \u1_m0_wo0_mtree_add4_0_o[9]~17_cout ;
wire \u1_m0_wo0_mtree_add4_0_o[9]~19_cout ;
wire \u1_m0_wo0_mtree_add4_0_o[9]~21_cout ;
wire \u1_m0_wo0_mtree_add4_0_o[9]~23_cout ;
wire \u1_m0_wo0_mtree_add4_0_o[9]~25_cout ;
wire \u1_m0_wo0_mtree_add4_0_o[9]~27_cout ;
wire \u1_m0_wo0_mtree_add4_0_o[9]~29_cout ;
wire \u1_m0_wo0_mtree_add4_0_o[9]~30_combout ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[1]~13 ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[2]~15 ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[3]~17 ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[4]~19 ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[5]~21 ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[6]~23 ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[7]~25 ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[8]~27 ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[9]~28_combout ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[8]~26_combout ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[7]~24_combout ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[6]~22_combout ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[5]~20_combout ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[4]~18_combout ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[3]~16_combout ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[2]~14_combout ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[1]~12_combout ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[0]~q ;
wire \u0_m0_wo0_mtree_add1_1_o[0]~15 ;
wire \u0_m0_wo0_mtree_add1_1_o[1]~17 ;
wire \u0_m0_wo0_mtree_add1_1_o[2]~19 ;
wire \u0_m0_wo0_mtree_add1_1_o[3]~21 ;
wire \u0_m0_wo0_mtree_add1_1_o[4]~23 ;
wire \u0_m0_wo0_mtree_add1_1_o[5]~25 ;
wire \u0_m0_wo0_mtree_add1_1_o[6]~27 ;
wire \u0_m0_wo0_mtree_add1_1_o[7]~29 ;
wire \u0_m0_wo0_mtree_add1_1_o[8]~31 ;
wire \u0_m0_wo0_mtree_add1_1_o[9]~32_combout ;
wire \u0_m0_wo0_mtree_add1_1_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[2]~14 ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[3]~16 ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[4]~18 ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[5]~20 ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[6]~22 ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[7]~24 ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[8]~26 ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[9]~27_combout ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[1]~14 ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[2]~16 ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[3]~18 ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[4]~20 ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[5]~22 ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[6]~24 ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[7]~26 ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[8]~27_combout ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[8]~25_combout ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[7]~25_combout ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[7]~23_combout ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[6]~23_combout ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[6]~21_combout ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[5]~21_combout ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[5]~19_combout ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[4]~19_combout ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[4]~17_combout ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[3]~17_combout ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[3]~15_combout ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[2]~15_combout ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[2]~13_combout ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[1]~13_combout ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[0]~q ;
wire \u0_m0_wo0_mtree_add0_4_o[1]~16 ;
wire \u0_m0_wo0_mtree_add0_4_o[2]~18 ;
wire \u0_m0_wo0_mtree_add0_4_o[3]~20 ;
wire \u0_m0_wo0_mtree_add0_4_o[4]~22 ;
wire \u0_m0_wo0_mtree_add0_4_o[5]~24 ;
wire \u0_m0_wo0_mtree_add0_4_o[6]~26 ;
wire \u0_m0_wo0_mtree_add0_4_o[7]~28 ;
wire \u0_m0_wo0_mtree_add0_4_o[8]~30 ;
wire \u0_m0_wo0_mtree_add0_4_o[9]~31_combout ;
wire \u0_m0_wo0_mtree_add0_4_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[1]~13 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[2]~15 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[3]~17 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[4]~19 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[5]~21 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[6]~23 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[7]~25 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[8]~27 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[9]~28_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[8]~26_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[7]~24_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[6]~22_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[5]~20_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[4]~18_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[3]~16_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[0]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[2]~14_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[2]~14 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[3]~16 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[4]~18 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[5]~20 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[6]~22 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[7]~24 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[8]~26 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[9]~27_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[9]~q ;
wire \u0_m0_wo0_mtree_add0_4_o[8]~29_combout ;
wire \u0_m0_wo0_mtree_add0_4_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[8]~25_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[8]~q ;
wire \u0_m0_wo0_mtree_add0_4_o[7]~27_combout ;
wire \u0_m0_wo0_mtree_add0_4_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[7]~23_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[7]~q ;
wire \u0_m0_wo0_mtree_add0_4_o[6]~25_combout ;
wire \u0_m0_wo0_mtree_add0_4_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[6]~21_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[6]~q ;
wire \u0_m0_wo0_mtree_add0_4_o[5]~23_combout ;
wire \u0_m0_wo0_mtree_add0_4_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[5]~19_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[5]~q ;
wire \u0_m0_wo0_mtree_add0_4_o[4]~21_combout ;
wire \u0_m0_wo0_mtree_add0_4_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[4]~17_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[4]~q ;
wire \u0_m0_wo0_mtree_add0_4_o[3]~19_combout ;
wire \u0_m0_wo0_mtree_add0_4_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[3]~15_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[3]~q ;
wire \u0_m0_wo0_mtree_add0_4_o[2]~17_combout ;
wire \u0_m0_wo0_mtree_add0_4_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[2]~13_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[2]~q ;
wire \u0_m0_wo0_mtree_add0_4_o[1]~15_combout ;
wire \u0_m0_wo0_mtree_add0_4_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[1]~12_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[0]~q ;
wire \u0_m0_wo0_mtree_add0_4_o[0]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[0]~q ;
wire \u0_m0_wo0_mtree_add1_2_o[0]~18 ;
wire \u0_m0_wo0_mtree_add1_2_o[1]~20 ;
wire \u0_m0_wo0_mtree_add1_2_o[2]~22 ;
wire \u0_m0_wo0_mtree_add1_2_o[3]~24 ;
wire \u0_m0_wo0_mtree_add1_2_o[4]~26 ;
wire \u0_m0_wo0_mtree_add1_2_o[5]~28 ;
wire \u0_m0_wo0_mtree_add1_2_o[6]~30 ;
wire \u0_m0_wo0_mtree_add1_2_o[7]~32 ;
wire \u0_m0_wo0_mtree_add1_2_o[8]~34 ;
wire \u0_m0_wo0_mtree_add1_2_o[9]~35_combout ;
wire \u0_m0_wo0_mtree_add1_2_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[1]~14 ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[2]~16 ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[3]~18 ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[4]~20 ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[5]~22 ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[6]~24 ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[7]~26 ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[8]~28 ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[9]~29_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[8]~27_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[7]~25_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[6]~23_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[5]~21_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[4]~19_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[0]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[3]~17_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[3]~14 ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[4]~16 ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[5]~18 ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[6]~20 ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[7]~22 ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[8]~24 ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[9]~25_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[1]~16 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[2]~18 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[3]~20 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[4]~22 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[5]~24 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[6]~26 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[7]~28 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[8]~30 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[9]~31_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[8]~29_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[7]~27_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[6]~25_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[0]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[5]~23_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[5]~14 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[6]~16 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[7]~18 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[8]~20 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[9]~21_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[8]~23_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[8]~19_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[7]~21_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[7]~17_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[6]~19_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[6]~15_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[5]~17_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[5]~13_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[4]~15_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[4]~21_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[3]~13_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[3]~19_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[2]~15_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[2]~17_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[1]~13_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[1]~15_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[0]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[0]~q ;
wire \u0_m0_wo0_mtree_add0_6_o[0]~20 ;
wire \u0_m0_wo0_mtree_add0_6_o[1]~22 ;
wire \u0_m0_wo0_mtree_add0_6_o[2]~24 ;
wire \u0_m0_wo0_mtree_add0_6_o[3]~26 ;
wire \u0_m0_wo0_mtree_add0_6_o[4]~28 ;
wire \u0_m0_wo0_mtree_add0_6_o[5]~30 ;
wire \u0_m0_wo0_mtree_add0_6_o[6]~32 ;
wire \u0_m0_wo0_mtree_add0_6_o[7]~34 ;
wire \u0_m0_wo0_mtree_add0_6_o[8]~36 ;
wire \u0_m0_wo0_mtree_add0_6_o[9]~37_combout ;
wire \u0_m0_wo0_mtree_add0_6_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[2]~14 ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[3]~16 ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[4]~18 ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[5]~20 ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[6]~22 ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[7]~24 ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[8]~26 ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[9]~27_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[8]~25_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[7]~23_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[6]~21_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[0]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[5]~19_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[5]~14 ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[6]~16 ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[7]~18 ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[8]~20 ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[9]~21_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[1]~20 ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[2]~22 ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[3]~24 ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[4]~26 ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[5]~28 ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[6]~30 ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[7]~32 ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[8]~34 ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[9]~35_combout ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[8]~19_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[8]~33_combout ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[7]~17_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[7]~31_combout ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[6]~15_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[6]~29_combout ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[5]~13_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[5]~27_combout ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[4]~17_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[4]~25_combout ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[3]~15_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[3]~23_combout ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[2]~13_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[2]~21_combout ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[1]~19_combout ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[0]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[0]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[0]~22 ;
wire \u0_m0_wo0_mtree_add0_7_o[1]~24 ;
wire \u0_m0_wo0_mtree_add0_7_o[2]~26 ;
wire \u0_m0_wo0_mtree_add0_7_o[3]~28 ;
wire \u0_m0_wo0_mtree_add0_7_o[4]~30 ;
wire \u0_m0_wo0_mtree_add0_7_o[5]~32 ;
wire \u0_m0_wo0_mtree_add0_7_o[6]~34 ;
wire \u0_m0_wo0_mtree_add0_7_o[7]~36 ;
wire \u0_m0_wo0_mtree_add0_7_o[8]~38 ;
wire \u0_m0_wo0_mtree_add0_7_o[9]~39_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[9]~q ;
wire \u0_m0_wo0_mtree_add0_6_o[8]~35_combout ;
wire \u0_m0_wo0_mtree_add0_6_o[8]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[8]~37_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[8]~q ;
wire \u0_m0_wo0_mtree_add0_6_o[7]~33_combout ;
wire \u0_m0_wo0_mtree_add0_6_o[7]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[7]~35_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[7]~q ;
wire \u0_m0_wo0_mtree_add0_6_o[6]~31_combout ;
wire \u0_m0_wo0_mtree_add0_6_o[6]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[6]~33_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[6]~q ;
wire \u0_m0_wo0_mtree_add0_6_o[5]~29_combout ;
wire \u0_m0_wo0_mtree_add0_6_o[5]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[5]~31_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[5]~q ;
wire \u0_m0_wo0_mtree_add0_6_o[4]~27_combout ;
wire \u0_m0_wo0_mtree_add0_6_o[4]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[4]~29_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[4]~q ;
wire \u0_m0_wo0_mtree_add0_6_o[3]~25_combout ;
wire \u0_m0_wo0_mtree_add0_6_o[3]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[3]~27_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[3]~q ;
wire \u0_m0_wo0_mtree_add0_6_o[2]~23_combout ;
wire \u0_m0_wo0_mtree_add0_6_o[2]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[2]~25_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[2]~q ;
wire \u0_m0_wo0_mtree_add0_6_o[1]~21_combout ;
wire \u0_m0_wo0_mtree_add0_6_o[1]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[1]~23_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[1]~q ;
wire \u0_m0_wo0_mtree_add0_6_o[0]~19_combout ;
wire \u0_m0_wo0_mtree_add0_6_o[0]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[0]~21_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[0]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[0]~22 ;
wire \u0_m0_wo0_mtree_add1_3_o[1]~24 ;
wire \u0_m0_wo0_mtree_add1_3_o[2]~26 ;
wire \u0_m0_wo0_mtree_add1_3_o[3]~28 ;
wire \u0_m0_wo0_mtree_add1_3_o[4]~30 ;
wire \u0_m0_wo0_mtree_add1_3_o[5]~32 ;
wire \u0_m0_wo0_mtree_add1_3_o[6]~34 ;
wire \u0_m0_wo0_mtree_add1_3_o[7]~36 ;
wire \u0_m0_wo0_mtree_add1_3_o[8]~38 ;
wire \u0_m0_wo0_mtree_add1_3_o[9]~39_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[9]~q ;
wire \u0_m0_wo0_mtree_add1_2_o[8]~33_combout ;
wire \u0_m0_wo0_mtree_add1_2_o[8]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[8]~37_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[8]~q ;
wire \u0_m0_wo0_mtree_add1_2_o[7]~31_combout ;
wire \u0_m0_wo0_mtree_add1_2_o[7]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[7]~35_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[7]~q ;
wire \u0_m0_wo0_mtree_add1_2_o[6]~29_combout ;
wire \u0_m0_wo0_mtree_add1_2_o[6]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[6]~33_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[6]~q ;
wire \u0_m0_wo0_mtree_add1_2_o[5]~27_combout ;
wire \u0_m0_wo0_mtree_add1_2_o[5]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[5]~31_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[5]~q ;
wire \u0_m0_wo0_mtree_add1_2_o[4]~25_combout ;
wire \u0_m0_wo0_mtree_add1_2_o[4]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[4]~29_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[4]~q ;
wire \u0_m0_wo0_mtree_add1_2_o[3]~23_combout ;
wire \u0_m0_wo0_mtree_add1_2_o[3]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[3]~27_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[3]~q ;
wire \u0_m0_wo0_mtree_add1_2_o[2]~21_combout ;
wire \u0_m0_wo0_mtree_add1_2_o[2]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[2]~25_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[2]~q ;
wire \u0_m0_wo0_mtree_add1_2_o[1]~19_combout ;
wire \u0_m0_wo0_mtree_add1_2_o[1]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[1]~23_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[1]~q ;
wire \u0_m0_wo0_mtree_add1_2_o[0]~17_combout ;
wire \u0_m0_wo0_mtree_add1_2_o[0]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[0]~21_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[0]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[0]~22 ;
wire \u0_m0_wo0_mtree_add2_1_o[1]~24 ;
wire \u0_m0_wo0_mtree_add2_1_o[2]~26 ;
wire \u0_m0_wo0_mtree_add2_1_o[3]~28 ;
wire \u0_m0_wo0_mtree_add2_1_o[4]~30 ;
wire \u0_m0_wo0_mtree_add2_1_o[5]~32 ;
wire \u0_m0_wo0_mtree_add2_1_o[6]~34 ;
wire \u0_m0_wo0_mtree_add2_1_o[7]~36 ;
wire \u0_m0_wo0_mtree_add2_1_o[8]~38 ;
wire \u0_m0_wo0_mtree_add2_1_o[9]~39_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[9]~q ;
wire \u0_m0_wo0_mtree_add1_1_o[8]~30_combout ;
wire \u0_m0_wo0_mtree_add1_1_o[8]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[8]~37_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[8]~q ;
wire \u0_m0_wo0_mtree_add1_1_o[7]~28_combout ;
wire \u0_m0_wo0_mtree_add1_1_o[7]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[7]~35_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[7]~q ;
wire \u0_m0_wo0_mtree_add1_1_o[6]~26_combout ;
wire \u0_m0_wo0_mtree_add1_1_o[6]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[6]~33_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[6]~q ;
wire \u0_m0_wo0_mtree_add1_1_o[5]~24_combout ;
wire \u0_m0_wo0_mtree_add1_1_o[5]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[5]~31_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[5]~q ;
wire \u0_m0_wo0_mtree_add1_1_o[4]~22_combout ;
wire \u0_m0_wo0_mtree_add1_1_o[4]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[4]~29_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[4]~q ;
wire \u0_m0_wo0_mtree_add1_1_o[3]~20_combout ;
wire \u0_m0_wo0_mtree_add1_1_o[3]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[3]~27_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[3]~q ;
wire \u0_m0_wo0_mtree_add1_1_o[2]~18_combout ;
wire \u0_m0_wo0_mtree_add1_1_o[2]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[2]~25_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[2]~q ;
wire \u0_m0_wo0_mtree_add1_1_o[1]~16_combout ;
wire \u0_m0_wo0_mtree_add1_1_o[1]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[1]~23_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[1]~q ;
wire \u0_m0_wo0_mtree_add1_1_o[0]~14_combout ;
wire \u0_m0_wo0_mtree_add1_1_o[0]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[0]~21_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[0]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[0]~22 ;
wire \u0_m0_wo0_mtree_add3_0_o[1]~24 ;
wire \u0_m0_wo0_mtree_add3_0_o[2]~26 ;
wire \u0_m0_wo0_mtree_add3_0_o[3]~28 ;
wire \u0_m0_wo0_mtree_add3_0_o[4]~30 ;
wire \u0_m0_wo0_mtree_add3_0_o[5]~32 ;
wire \u0_m0_wo0_mtree_add3_0_o[6]~34 ;
wire \u0_m0_wo0_mtree_add3_0_o[7]~36 ;
wire \u0_m0_wo0_mtree_add3_0_o[8]~38 ;
wire \u0_m0_wo0_mtree_add3_0_o[9]~39_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[2]~14 ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[3]~16 ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[4]~18 ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[5]~20 ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[6]~22 ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[7]~24 ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[8]~26 ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[9]~27_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[8]~25_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[7]~23_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[6]~21_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[0]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[5]~19_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[5]~14 ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[6]~16 ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[7]~18 ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[8]~20 ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[9]~21_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[1]~16 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[2]~18 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[3]~20 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[4]~22 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[5]~24 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[6]~26 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[7]~28 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[8]~30 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[9]~31_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[8]~29_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[7]~27_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[6]~25_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[0]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[5]~23_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[5]~14 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[6]~16 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[7]~18 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[8]~20 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[9]~21_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[8]~19_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[8]~19_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[7]~17_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[7]~17_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[6]~15_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[6]~15_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[5]~13_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[5]~13_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[4]~17_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[4]~21_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[3]~15_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[3]~19_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[2]~13_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[2]~17_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[1]~15_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[0]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[0]~q ;
wire \u0_m0_wo0_mtree_add0_8_o[0]~20 ;
wire \u0_m0_wo0_mtree_add0_8_o[1]~22 ;
wire \u0_m0_wo0_mtree_add0_8_o[2]~24 ;
wire \u0_m0_wo0_mtree_add0_8_o[3]~26 ;
wire \u0_m0_wo0_mtree_add0_8_o[4]~28 ;
wire \u0_m0_wo0_mtree_add0_8_o[5]~30 ;
wire \u0_m0_wo0_mtree_add0_8_o[6]~32 ;
wire \u0_m0_wo0_mtree_add0_8_o[7]~34 ;
wire \u0_m0_wo0_mtree_add0_8_o[8]~36 ;
wire \u0_m0_wo0_mtree_add0_8_o[9]~37_combout ;
wire \u0_m0_wo0_mtree_add0_8_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[1]~14 ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[2]~16 ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[3]~18 ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[4]~20 ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[5]~22 ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[6]~24 ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[7]~26 ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[8]~28 ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[9]~29_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[8]~27_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[7]~25_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[6]~23_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[5]~21_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[4]~19_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[0]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[3]~17_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[3]~14 ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[4]~16 ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[5]~18 ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[6]~20 ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[7]~22 ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[8]~24 ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[9]~25_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[9]~q ;
wire \u0_m0_wo0_mtree_add0_8_o[8]~35_combout ;
wire \u0_m0_wo0_mtree_add0_8_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[8]~23_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[8]~q ;
wire \u0_m0_wo0_mtree_add0_8_o[7]~33_combout ;
wire \u0_m0_wo0_mtree_add0_8_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[7]~21_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[7]~q ;
wire \u0_m0_wo0_mtree_add0_8_o[6]~31_combout ;
wire \u0_m0_wo0_mtree_add0_8_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[6]~19_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[6]~q ;
wire \u0_m0_wo0_mtree_add0_8_o[5]~29_combout ;
wire \u0_m0_wo0_mtree_add0_8_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[5]~17_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[5]~q ;
wire \u0_m0_wo0_mtree_add0_8_o[4]~27_combout ;
wire \u0_m0_wo0_mtree_add0_8_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[4]~15_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[4]~q ;
wire \u0_m0_wo0_mtree_add0_8_o[3]~25_combout ;
wire \u0_m0_wo0_mtree_add0_8_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[3]~13_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[3]~q ;
wire \u0_m0_wo0_mtree_add0_8_o[2]~23_combout ;
wire \u0_m0_wo0_mtree_add0_8_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[2]~15_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[2]~q ;
wire \u0_m0_wo0_mtree_add0_8_o[1]~21_combout ;
wire \u0_m0_wo0_mtree_add0_8_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[1]~13_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[1]~q ;
wire \u0_m0_wo0_mtree_add0_8_o[0]~19_combout ;
wire \u0_m0_wo0_mtree_add0_8_o[0]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[0]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[0]~21 ;
wire \u0_m0_wo0_mtree_add1_4_o[1]~23 ;
wire \u0_m0_wo0_mtree_add1_4_o[2]~25 ;
wire \u0_m0_wo0_mtree_add1_4_o[3]~27 ;
wire \u0_m0_wo0_mtree_add1_4_o[4]~29 ;
wire \u0_m0_wo0_mtree_add1_4_o[5]~31 ;
wire \u0_m0_wo0_mtree_add1_4_o[6]~33 ;
wire \u0_m0_wo0_mtree_add1_4_o[7]~35 ;
wire \u0_m0_wo0_mtree_add1_4_o[8]~37 ;
wire \u0_m0_wo0_mtree_add1_4_o[9]~38_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[1]~13 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[2]~15 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[3]~17 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[4]~19 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[5]~21 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[6]~23 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[7]~25 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[8]~27 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[9]~28_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[8]~26_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[7]~24_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[6]~22_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[5]~20_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[4]~18_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[3]~16_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[0]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[2]~14_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[2]~14 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[3]~16 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[4]~18 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[5]~20 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[6]~22 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[7]~24 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[8]~26 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[9]~27_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[1]~14 ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[2]~16 ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[3]~18 ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[4]~20 ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[5]~22 ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[6]~24 ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[7]~26 ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[8]~27_combout ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[8]~25_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[7]~25_combout ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[7]~23_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[6]~23_combout ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[6]~21_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[5]~21_combout ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[5]~19_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[4]~19_combout ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[4]~17_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[3]~17_combout ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[3]~15_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[2]~15_combout ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[2]~13_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[1]~13_combout ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[1]~12_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[0]~q ;
wire \u0_m0_wo0_mtree_add0_10_o[1]~16 ;
wire \u0_m0_wo0_mtree_add0_10_o[2]~18 ;
wire \u0_m0_wo0_mtree_add0_10_o[3]~20 ;
wire \u0_m0_wo0_mtree_add0_10_o[4]~22 ;
wire \u0_m0_wo0_mtree_add0_10_o[5]~24 ;
wire \u0_m0_wo0_mtree_add0_10_o[6]~26 ;
wire \u0_m0_wo0_mtree_add0_10_o[7]~28 ;
wire \u0_m0_wo0_mtree_add0_10_o[8]~30 ;
wire \u0_m0_wo0_mtree_add0_10_o[9]~31_combout ;
wire \u0_m0_wo0_mtree_add0_10_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[2]~14 ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[3]~16 ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[4]~18 ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[5]~20 ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[6]~22 ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[7]~24 ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[8]~26 ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[9]~27_combout ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[9]~q ;
wire \u0_m0_wo0_mtree_add0_10_o[8]~29_combout ;
wire \u0_m0_wo0_mtree_add0_10_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[8]~25_combout ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[8]~q ;
wire \u0_m0_wo0_mtree_add0_10_o[7]~27_combout ;
wire \u0_m0_wo0_mtree_add0_10_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[7]~23_combout ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[7]~q ;
wire \u0_m0_wo0_mtree_add0_10_o[6]~25_combout ;
wire \u0_m0_wo0_mtree_add0_10_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[6]~21_combout ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[6]~q ;
wire \u0_m0_wo0_mtree_add0_10_o[5]~23_combout ;
wire \u0_m0_wo0_mtree_add0_10_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[5]~19_combout ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[5]~q ;
wire \u0_m0_wo0_mtree_add0_10_o[4]~21_combout ;
wire \u0_m0_wo0_mtree_add0_10_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[4]~17_combout ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[4]~q ;
wire \u0_m0_wo0_mtree_add0_10_o[3]~19_combout ;
wire \u0_m0_wo0_mtree_add0_10_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[3]~15_combout ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[3]~q ;
wire \u0_m0_wo0_mtree_add0_10_o[2]~17_combout ;
wire \u0_m0_wo0_mtree_add0_10_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[2]~13_combout ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[2]~q ;
wire \u0_m0_wo0_mtree_add0_10_o[1]~15_combout ;
wire \u0_m0_wo0_mtree_add0_10_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[0]~q ;
wire \u0_m0_wo0_mtree_add0_10_o[0]~q ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[0]~q ;
wire \u0_m0_wo0_mtree_add1_5_o[0]~18 ;
wire \u0_m0_wo0_mtree_add1_5_o[1]~20 ;
wire \u0_m0_wo0_mtree_add1_5_o[2]~22 ;
wire \u0_m0_wo0_mtree_add1_5_o[3]~24 ;
wire \u0_m0_wo0_mtree_add1_5_o[4]~26 ;
wire \u0_m0_wo0_mtree_add1_5_o[5]~28 ;
wire \u0_m0_wo0_mtree_add1_5_o[6]~30 ;
wire \u0_m0_wo0_mtree_add1_5_o[7]~32 ;
wire \u0_m0_wo0_mtree_add1_5_o[8]~34 ;
wire \u0_m0_wo0_mtree_add1_5_o[9]~35_combout ;
wire \u0_m0_wo0_mtree_add1_5_o[9]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[8]~36_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[8]~q ;
wire \u0_m0_wo0_mtree_add1_5_o[8]~33_combout ;
wire \u0_m0_wo0_mtree_add1_5_o[8]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[7]~34_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[7]~q ;
wire \u0_m0_wo0_mtree_add1_5_o[7]~31_combout ;
wire \u0_m0_wo0_mtree_add1_5_o[7]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[6]~32_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[6]~q ;
wire \u0_m0_wo0_mtree_add1_5_o[6]~29_combout ;
wire \u0_m0_wo0_mtree_add1_5_o[6]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[5]~30_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[5]~q ;
wire \u0_m0_wo0_mtree_add1_5_o[5]~27_combout ;
wire \u0_m0_wo0_mtree_add1_5_o[5]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[4]~28_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[4]~q ;
wire \u0_m0_wo0_mtree_add1_5_o[4]~25_combout ;
wire \u0_m0_wo0_mtree_add1_5_o[4]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[3]~26_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[3]~q ;
wire \u0_m0_wo0_mtree_add1_5_o[3]~23_combout ;
wire \u0_m0_wo0_mtree_add1_5_o[3]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[2]~24_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[2]~q ;
wire \u0_m0_wo0_mtree_add1_5_o[2]~21_combout ;
wire \u0_m0_wo0_mtree_add1_5_o[2]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[1]~22_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[1]~q ;
wire \u0_m0_wo0_mtree_add1_5_o[1]~19_combout ;
wire \u0_m0_wo0_mtree_add1_5_o[1]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[0]~20_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[0]~q ;
wire \u0_m0_wo0_mtree_add1_5_o[0]~17_combout ;
wire \u0_m0_wo0_mtree_add1_5_o[0]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[0]~22 ;
wire \u0_m0_wo0_mtree_add2_2_o[1]~24 ;
wire \u0_m0_wo0_mtree_add2_2_o[2]~26 ;
wire \u0_m0_wo0_mtree_add2_2_o[3]~28 ;
wire \u0_m0_wo0_mtree_add2_2_o[4]~30 ;
wire \u0_m0_wo0_mtree_add2_2_o[5]~32 ;
wire \u0_m0_wo0_mtree_add2_2_o[6]~34 ;
wire \u0_m0_wo0_mtree_add2_2_o[7]~36 ;
wire \u0_m0_wo0_mtree_add2_2_o[8]~38 ;
wire \u0_m0_wo0_mtree_add2_2_o[9]~39_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[1]~13 ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[2]~15 ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[3]~17 ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[4]~19 ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[5]~21 ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[6]~23 ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[7]~25 ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[8]~27 ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[9]~28_combout ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[9]~q ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[8]~26_combout ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[8]~q ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[7]~24_combout ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[7]~q ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[6]~22_combout ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[6]~q ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[5]~20_combout ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[5]~q ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[4]~18_combout ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[4]~q ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[3]~16_combout ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[3]~q ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[2]~14_combout ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[2]~q ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[1]~12_combout ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[1]~q ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[0]~q ;
wire \u0_m0_wo0_mtree_add0_12_o[0]~15 ;
wire \u0_m0_wo0_mtree_add0_12_o[1]~17 ;
wire \u0_m0_wo0_mtree_add0_12_o[2]~19 ;
wire \u0_m0_wo0_mtree_add0_12_o[3]~21 ;
wire \u0_m0_wo0_mtree_add0_12_o[4]~23 ;
wire \u0_m0_wo0_mtree_add0_12_o[5]~25 ;
wire \u0_m0_wo0_mtree_add0_12_o[6]~27 ;
wire \u0_m0_wo0_mtree_add0_12_o[7]~29 ;
wire \u0_m0_wo0_mtree_add0_12_o[8]~31 ;
wire \u0_m0_wo0_mtree_add0_12_o[9]~32_combout ;
wire \u0_m0_wo0_mtree_add0_12_o[9]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[8]~37_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[8]~q ;
wire \u0_m0_wo0_mtree_add0_12_o[8]~30_combout ;
wire \u0_m0_wo0_mtree_add0_12_o[8]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[7]~35_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[7]~q ;
wire \u0_m0_wo0_mtree_add0_12_o[7]~28_combout ;
wire \u0_m0_wo0_mtree_add0_12_o[7]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[6]~33_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[6]~q ;
wire \u0_m0_wo0_mtree_add0_12_o[6]~26_combout ;
wire \u0_m0_wo0_mtree_add0_12_o[6]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[5]~31_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[5]~q ;
wire \u0_m0_wo0_mtree_add0_12_o[5]~24_combout ;
wire \u0_m0_wo0_mtree_add0_12_o[5]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[4]~29_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[4]~q ;
wire \u0_m0_wo0_mtree_add0_12_o[4]~22_combout ;
wire \u0_m0_wo0_mtree_add0_12_o[4]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[3]~27_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[3]~q ;
wire \u0_m0_wo0_mtree_add0_12_o[3]~20_combout ;
wire \u0_m0_wo0_mtree_add0_12_o[3]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[2]~25_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[2]~q ;
wire \u0_m0_wo0_mtree_add0_12_o[2]~18_combout ;
wire \u0_m0_wo0_mtree_add0_12_o[2]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[1]~23_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[1]~q ;
wire \u0_m0_wo0_mtree_add0_12_o[1]~16_combout ;
wire \u0_m0_wo0_mtree_add0_12_o[1]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[0]~21_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[0]~q ;
wire \u0_m0_wo0_mtree_add0_12_o[0]~14_combout ;
wire \u0_m0_wo0_mtree_add0_12_o[0]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[0]~22 ;
wire \u0_m0_wo0_mtree_add3_1_o[1]~24 ;
wire \u0_m0_wo0_mtree_add3_1_o[2]~26 ;
wire \u0_m0_wo0_mtree_add3_1_o[3]~28 ;
wire \u0_m0_wo0_mtree_add3_1_o[4]~30 ;
wire \u0_m0_wo0_mtree_add3_1_o[5]~32 ;
wire \u0_m0_wo0_mtree_add3_1_o[6]~34 ;
wire \u0_m0_wo0_mtree_add3_1_o[7]~36 ;
wire \u0_m0_wo0_mtree_add3_1_o[8]~38 ;
wire \u0_m0_wo0_mtree_add3_1_o[9]~39_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[9]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[8]~37_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[8]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[8]~37_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[8]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[7]~35_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[7]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[7]~35_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[7]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[6]~33_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[6]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[6]~33_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[6]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[5]~31_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[5]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[5]~31_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[5]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[4]~29_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[4]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[4]~29_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[4]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[3]~27_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[3]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[3]~27_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[3]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[2]~25_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[2]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[2]~25_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[2]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[1]~23_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[1]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[1]~23_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[1]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[0]~21_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[0]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[0]~21_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[0]~q ;
wire \u0_m0_wo0_mtree_add4_0_o[9]~13_cout ;
wire \u0_m0_wo0_mtree_add4_0_o[9]~15_cout ;
wire \u0_m0_wo0_mtree_add4_0_o[9]~17_cout ;
wire \u0_m0_wo0_mtree_add4_0_o[9]~19_cout ;
wire \u0_m0_wo0_mtree_add4_0_o[9]~21_cout ;
wire \u0_m0_wo0_mtree_add4_0_o[9]~23_cout ;
wire \u0_m0_wo0_mtree_add4_0_o[9]~25_cout ;
wire \u0_m0_wo0_mtree_add4_0_o[9]~27_cout ;
wire \u0_m0_wo0_mtree_add4_0_o[9]~29_cout ;
wire \u0_m0_wo0_mtree_add4_0_o[9]~30_combout ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[9]~29 ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[10]~31 ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[11]~33 ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[12]~34_combout ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[11]~32_combout ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[10]~30_combout ;
wire \u0_m0_wo0_mtree_mult1_5_sub_0_o[10]~q ;
wire \u0_m0_wo0_mtree_add1_1_o[9]~33 ;
wire \u0_m0_wo0_mtree_add1_1_o[10]~35 ;
wire \u0_m0_wo0_mtree_add1_1_o[11]~37 ;
wire \u0_m0_wo0_mtree_add1_1_o[12]~39 ;
wire \u0_m0_wo0_mtree_add1_1_o[15]~40_combout ;
wire \u0_m0_wo0_mtree_add1_1_o[15]~q ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[9]~28 ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[10]~30 ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[11]~32 ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[12]~34 ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[13]~36 ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[14]~37_combout ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[14]~q ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[8]~28 ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[9]~30 ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[10]~32 ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[11]~34 ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[12]~36 ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[13]~37_combout ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[13]~q ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[13]~35_combout ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[13]~q ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[12]~35_combout ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[12]~33_combout ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[11]~33_combout ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[11]~31_combout ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[10]~31_combout ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[10]~q ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[10]~29_combout ;
wire \u0_m0_wo0_mtree_mult1_8_sub_1_o[10]~q ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[9]~29_combout ;
wire \u0_m0_wo0_mtree_mult1_9_add_1_o[9]~q ;
wire \u0_m0_wo0_mtree_add0_4_o[9]~32 ;
wire \u0_m0_wo0_mtree_add0_4_o[10]~34 ;
wire \u0_m0_wo0_mtree_add0_4_o[11]~36 ;
wire \u0_m0_wo0_mtree_add0_4_o[12]~38 ;
wire \u0_m0_wo0_mtree_add0_4_o[13]~40 ;
wire \u0_m0_wo0_mtree_add0_4_o[14]~42 ;
wire \u0_m0_wo0_mtree_add0_4_o[15]~43_combout ;
wire \u0_m0_wo0_mtree_add0_4_o[15]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[9]~29 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[10]~31 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[11]~33 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[12]~34_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[11]~32_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[10]~30_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_0_o[10]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[9]~28 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[10]~30 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[11]~32 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[12]~34 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[13]~36 ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[14]~37_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[14]~q ;
wire \u0_m0_wo0_mtree_add0_4_o[14]~41_combout ;
wire \u0_m0_wo0_mtree_add0_4_o[14]~q ;
wire \u0_m0_wo0_mtree_add0_4_o[13]~39_combout ;
wire \u0_m0_wo0_mtree_add0_4_o[13]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[13]~35_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[13]~q ;
wire \u0_m0_wo0_mtree_add0_4_o[12]~37_combout ;
wire \u0_m0_wo0_mtree_add0_4_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[12]~33_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[12]~q ;
wire \u0_m0_wo0_mtree_add0_4_o[11]~35_combout ;
wire \u0_m0_wo0_mtree_add0_4_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[11]~31_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[11]~q ;
wire \u0_m0_wo0_mtree_add0_4_o[10]~33_combout ;
wire \u0_m0_wo0_mtree_add0_4_o[10]~q ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[10]~29_combout ;
wire \u0_m0_wo0_mtree_mult1_10_sub_2_o[10]~q ;
wire \u0_m0_wo0_mtree_add1_2_o[9]~36 ;
wire \u0_m0_wo0_mtree_add1_2_o[10]~38 ;
wire \u0_m0_wo0_mtree_add1_2_o[11]~40 ;
wire \u0_m0_wo0_mtree_add1_2_o[12]~42 ;
wire \u0_m0_wo0_mtree_add1_2_o[13]~44 ;
wire \u0_m0_wo0_mtree_add1_2_o[14]~46 ;
wire \u0_m0_wo0_mtree_add1_2_o[15]~48 ;
wire \u0_m0_wo0_mtree_add1_2_o[17]~49_combout ;
wire \u0_m0_wo0_mtree_add1_2_o[17]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[9]~30 ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[10]~32 ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[11]~34 ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[12]~36 ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[13]~37_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[13]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[12]~35_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[11]~33_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[10]~31_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_1_o[10]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[9]~26 ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[10]~28 ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[11]~30 ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[12]~32 ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[13]~34 ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[14]~36 ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[15]~37_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[15]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[9]~32 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[10]~34 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[11]~36 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[12]~38 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[13]~40 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[14]~42 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[15]~43_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[15]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[14]~41_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[14]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[13]~39_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[13]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[12]~37_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[11]~35_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[10]~33_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_1_o[10]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[9]~22 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[10]~24 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[11]~26 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[12]~28 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[13]~30 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[14]~32 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[15]~34 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[16]~36 ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[17]~37_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[17]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[16]~35_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[16]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[15]~33_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[15]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[14]~35_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[14]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[14]~31_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[14]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[13]~33_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[13]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[13]~29_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[13]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[12]~31_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[12]~27_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[11]~29_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[11]~25_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[10]~27_combout ;
wire \u0_m0_wo0_mtree_mult1_12_add_3_o[10]~q ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[10]~23_combout ;
wire \u0_m0_wo0_mtree_mult1_13_sub_3_o[10]~q ;
wire \u0_m0_wo0_mtree_add0_6_o[9]~38 ;
wire \u0_m0_wo0_mtree_add0_6_o[10]~40 ;
wire \u0_m0_wo0_mtree_add0_6_o[11]~42 ;
wire \u0_m0_wo0_mtree_add0_6_o[12]~44 ;
wire \u0_m0_wo0_mtree_add0_6_o[13]~46 ;
wire \u0_m0_wo0_mtree_add0_6_o[14]~48 ;
wire \u0_m0_wo0_mtree_add0_6_o[15]~50 ;
wire \u0_m0_wo0_mtree_add0_6_o[16]~52 ;
wire \u0_m0_wo0_mtree_add0_6_o[17]~54 ;
wire \u0_m0_wo0_mtree_add0_6_o[18]~55_combout ;
wire \u0_m0_wo0_mtree_add0_6_o[18]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[9]~28 ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[10]~30 ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[11]~32 ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[12]~34 ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[13]~36 ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[14]~37_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[14]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[13]~35_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[13]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[12]~33_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[11]~31_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[10]~29_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_1_o[10]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[9]~22 ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[10]~24 ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[11]~26 ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[12]~28 ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[13]~30 ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[14]~32 ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[15]~34 ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[16]~36 ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[17]~37_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[17]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[9]~36 ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[10]~38 ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[11]~40 ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[12]~42 ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[13]~44 ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[14]~46 ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[15]~48 ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[16]~50 ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[17]~52 ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[18]~54 ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[19]~55_combout ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[19]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[18]~53_combout ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[18]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[17]~51_combout ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[17]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[16]~35_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[16]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[16]~49_combout ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[16]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[15]~33_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[15]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[15]~47_combout ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[15]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[14]~31_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[14]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[14]~45_combout ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[14]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[13]~29_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[13]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[13]~43_combout ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[13]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[12]~27_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[12]~41_combout ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[11]~25_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[11]~39_combout ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[10]~23_combout ;
wire \u0_m0_wo0_mtree_mult1_14_add_3_o[10]~q ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[10]~37_combout ;
wire \u0_m0_wo0_mtree_mult1_15_sub_1_o[10]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[9]~40 ;
wire \u0_m0_wo0_mtree_add0_7_o[10]~42 ;
wire \u0_m0_wo0_mtree_add0_7_o[11]~44 ;
wire \u0_m0_wo0_mtree_add0_7_o[12]~46 ;
wire \u0_m0_wo0_mtree_add0_7_o[13]~48 ;
wire \u0_m0_wo0_mtree_add0_7_o[14]~50 ;
wire \u0_m0_wo0_mtree_add0_7_o[15]~52 ;
wire \u0_m0_wo0_mtree_add0_7_o[16]~54 ;
wire \u0_m0_wo0_mtree_add0_7_o[17]~56 ;
wire \u0_m0_wo0_mtree_add0_7_o[18]~58 ;
wire \u0_m0_wo0_mtree_add0_7_o[19]~60 ;
wire \u0_m0_wo0_mtree_add0_7_o[20]~61_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[20]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[19]~59_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[19]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[18]~57_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[18]~q ;
wire \u0_m0_wo0_mtree_add0_6_o[17]~53_combout ;
wire \u0_m0_wo0_mtree_add0_6_o[17]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[17]~55_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[17]~q ;
wire \u0_m0_wo0_mtree_add0_6_o[16]~51_combout ;
wire \u0_m0_wo0_mtree_add0_6_o[16]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[16]~53_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[16]~q ;
wire \u0_m0_wo0_mtree_add0_6_o[15]~49_combout ;
wire \u0_m0_wo0_mtree_add0_6_o[15]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[15]~51_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[15]~q ;
wire \u0_m0_wo0_mtree_add0_6_o[14]~47_combout ;
wire \u0_m0_wo0_mtree_add0_6_o[14]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[14]~49_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[14]~q ;
wire \u0_m0_wo0_mtree_add0_6_o[13]~45_combout ;
wire \u0_m0_wo0_mtree_add0_6_o[13]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[13]~47_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[13]~q ;
wire \u0_m0_wo0_mtree_add0_6_o[12]~43_combout ;
wire \u0_m0_wo0_mtree_add0_6_o[12]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[12]~45_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[12]~q ;
wire \u0_m0_wo0_mtree_add0_6_o[11]~41_combout ;
wire \u0_m0_wo0_mtree_add0_6_o[11]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[11]~43_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[11]~q ;
wire \u0_m0_wo0_mtree_add0_6_o[10]~39_combout ;
wire \u0_m0_wo0_mtree_add0_6_o[10]~q ;
wire \u0_m0_wo0_mtree_add0_7_o[10]~41_combout ;
wire \u0_m0_wo0_mtree_add0_7_o[10]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[9]~40 ;
wire \u0_m0_wo0_mtree_add1_3_o[10]~42 ;
wire \u0_m0_wo0_mtree_add1_3_o[11]~44 ;
wire \u0_m0_wo0_mtree_add1_3_o[12]~46 ;
wire \u0_m0_wo0_mtree_add1_3_o[13]~48 ;
wire \u0_m0_wo0_mtree_add1_3_o[14]~50 ;
wire \u0_m0_wo0_mtree_add1_3_o[15]~52 ;
wire \u0_m0_wo0_mtree_add1_3_o[16]~54 ;
wire \u0_m0_wo0_mtree_add1_3_o[17]~56 ;
wire \u0_m0_wo0_mtree_add1_3_o[18]~58 ;
wire \u0_m0_wo0_mtree_add1_3_o[19]~60 ;
wire \u0_m0_wo0_mtree_add1_3_o[20]~61_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[20]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[19]~59_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[19]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[18]~57_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[18]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[17]~55_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[17]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[16]~53_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[16]~q ;
wire \u0_m0_wo0_mtree_add1_2_o[15]~47_combout ;
wire \u0_m0_wo0_mtree_add1_2_o[15]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[15]~51_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[15]~q ;
wire \u0_m0_wo0_mtree_add1_2_o[14]~45_combout ;
wire \u0_m0_wo0_mtree_add1_2_o[14]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[14]~49_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[14]~q ;
wire \u0_m0_wo0_mtree_add1_2_o[13]~43_combout ;
wire \u0_m0_wo0_mtree_add1_2_o[13]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[13]~47_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[13]~q ;
wire \u0_m0_wo0_mtree_add1_2_o[12]~41_combout ;
wire \u0_m0_wo0_mtree_add1_2_o[12]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[12]~45_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[12]~q ;
wire \u0_m0_wo0_mtree_add1_2_o[11]~39_combout ;
wire \u0_m0_wo0_mtree_add1_2_o[11]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[11]~43_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[11]~q ;
wire \u0_m0_wo0_mtree_add1_2_o[10]~37_combout ;
wire \u0_m0_wo0_mtree_add1_2_o[10]~q ;
wire \u0_m0_wo0_mtree_add1_3_o[10]~41_combout ;
wire \u0_m0_wo0_mtree_add1_3_o[10]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[9]~40 ;
wire \u0_m0_wo0_mtree_add2_1_o[10]~42 ;
wire \u0_m0_wo0_mtree_add2_1_o[11]~44 ;
wire \u0_m0_wo0_mtree_add2_1_o[12]~46 ;
wire \u0_m0_wo0_mtree_add2_1_o[13]~48 ;
wire \u0_m0_wo0_mtree_add2_1_o[14]~50 ;
wire \u0_m0_wo0_mtree_add2_1_o[15]~52 ;
wire \u0_m0_wo0_mtree_add2_1_o[16]~54 ;
wire \u0_m0_wo0_mtree_add2_1_o[17]~56 ;
wire \u0_m0_wo0_mtree_add2_1_o[18]~58 ;
wire \u0_m0_wo0_mtree_add2_1_o[19]~60 ;
wire \u0_m0_wo0_mtree_add2_1_o[20]~61_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[20]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[19]~59_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[19]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[18]~57_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[18]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[17]~55_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[17]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[16]~53_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[16]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[15]~51_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[15]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[14]~49_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[14]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[13]~47_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[13]~q ;
wire \u0_m0_wo0_mtree_add1_1_o[12]~38_combout ;
wire \u0_m0_wo0_mtree_add1_1_o[12]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[12]~45_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[12]~q ;
wire \u0_m0_wo0_mtree_add1_1_o[11]~36_combout ;
wire \u0_m0_wo0_mtree_add1_1_o[11]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[11]~43_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[11]~q ;
wire \u0_m0_wo0_mtree_add1_1_o[10]~34_combout ;
wire \u0_m0_wo0_mtree_add1_1_o[10]~q ;
wire \u0_m0_wo0_mtree_add2_1_o[10]~41_combout ;
wire \u0_m0_wo0_mtree_add2_1_o[10]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[9]~40 ;
wire \u0_m0_wo0_mtree_add3_0_o[10]~42 ;
wire \u0_m0_wo0_mtree_add3_0_o[11]~44 ;
wire \u0_m0_wo0_mtree_add3_0_o[12]~46 ;
wire \u0_m0_wo0_mtree_add3_0_o[13]~48 ;
wire \u0_m0_wo0_mtree_add3_0_o[14]~50 ;
wire \u0_m0_wo0_mtree_add3_0_o[15]~52 ;
wire \u0_m0_wo0_mtree_add3_0_o[16]~54 ;
wire \u0_m0_wo0_mtree_add3_0_o[17]~56 ;
wire \u0_m0_wo0_mtree_add3_0_o[18]~58 ;
wire \u0_m0_wo0_mtree_add3_0_o[19]~60 ;
wire \u0_m0_wo0_mtree_add3_0_o[20]~61_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[20]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[9]~28 ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[10]~30 ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[11]~32 ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[12]~34 ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[13]~36 ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[14]~37_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[14]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[13]~35_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[13]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[12]~33_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[11]~31_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[10]~29_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_1_o[10]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[9]~22 ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[10]~24 ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[11]~26 ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[12]~28 ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[13]~30 ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[14]~32 ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[15]~34 ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[16]~36 ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[17]~37_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[17]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[9]~32 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[10]~34 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[11]~36 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[12]~38 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[13]~40 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[14]~42 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[15]~43_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[15]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[14]~41_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[14]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[13]~39_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[13]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[12]~37_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[11]~35_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[10]~33_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_1_o[10]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[9]~22 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[10]~24 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[11]~26 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[12]~28 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[13]~30 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[14]~32 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[15]~34 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[16]~36 ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[17]~37_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[17]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[16]~35_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[16]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[16]~35_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[16]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[15]~33_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[15]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[15]~33_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[15]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[14]~31_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[14]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[14]~31_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[14]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[13]~29_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[13]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[13]~29_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[13]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[12]~27_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[12]~27_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[11]~25_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[11]~25_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[10]~23_combout ;
wire \u0_m0_wo0_mtree_mult1_16_add_3_o[10]~q ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[10]~23_combout ;
wire \u0_m0_wo0_mtree_mult1_17_sub_3_o[10]~q ;
wire \u0_m0_wo0_mtree_add0_8_o[9]~38 ;
wire \u0_m0_wo0_mtree_add0_8_o[10]~40 ;
wire \u0_m0_wo0_mtree_add0_8_o[11]~42 ;
wire \u0_m0_wo0_mtree_add0_8_o[12]~44 ;
wire \u0_m0_wo0_mtree_add0_8_o[13]~46 ;
wire \u0_m0_wo0_mtree_add0_8_o[14]~48 ;
wire \u0_m0_wo0_mtree_add0_8_o[15]~50 ;
wire \u0_m0_wo0_mtree_add0_8_o[16]~52 ;
wire \u0_m0_wo0_mtree_add0_8_o[17]~54 ;
wire \u0_m0_wo0_mtree_add0_8_o[18]~55_combout ;
wire \u0_m0_wo0_mtree_add0_8_o[18]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[9]~30 ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[10]~32 ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[11]~34 ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[12]~36 ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[13]~37_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[13]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[12]~35_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[11]~33_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[10]~31_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_1_o[10]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[9]~26 ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[10]~28 ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[11]~30 ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[12]~32 ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[13]~34 ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[14]~36 ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[15]~37_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[15]~q ;
wire \u0_m0_wo0_mtree_add0_8_o[17]~53_combout ;
wire \u0_m0_wo0_mtree_add0_8_o[17]~q ;
wire \u0_m0_wo0_mtree_add0_8_o[16]~51_combout ;
wire \u0_m0_wo0_mtree_add0_8_o[16]~q ;
wire \u0_m0_wo0_mtree_add0_8_o[15]~49_combout ;
wire \u0_m0_wo0_mtree_add0_8_o[15]~q ;
wire \u0_m0_wo0_mtree_add0_8_o[14]~47_combout ;
wire \u0_m0_wo0_mtree_add0_8_o[14]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[14]~35_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[14]~q ;
wire \u0_m0_wo0_mtree_add0_8_o[13]~45_combout ;
wire \u0_m0_wo0_mtree_add0_8_o[13]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[13]~33_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[13]~q ;
wire \u0_m0_wo0_mtree_add0_8_o[12]~43_combout ;
wire \u0_m0_wo0_mtree_add0_8_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[12]~31_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[12]~q ;
wire \u0_m0_wo0_mtree_add0_8_o[11]~41_combout ;
wire \u0_m0_wo0_mtree_add0_8_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[11]~29_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[11]~q ;
wire \u0_m0_wo0_mtree_add0_8_o[10]~39_combout ;
wire \u0_m0_wo0_mtree_add0_8_o[10]~q ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[10]~27_combout ;
wire \u0_m0_wo0_mtree_mult1_18_add_3_o[10]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[9]~39 ;
wire \u0_m0_wo0_mtree_add1_4_o[10]~41 ;
wire \u0_m0_wo0_mtree_add1_4_o[11]~43 ;
wire \u0_m0_wo0_mtree_add1_4_o[12]~45 ;
wire \u0_m0_wo0_mtree_add1_4_o[13]~47 ;
wire \u0_m0_wo0_mtree_add1_4_o[14]~49 ;
wire \u0_m0_wo0_mtree_add1_4_o[15]~51 ;
wire \u0_m0_wo0_mtree_add1_4_o[16]~53 ;
wire \u0_m0_wo0_mtree_add1_4_o[17]~55 ;
wire \u0_m0_wo0_mtree_add1_4_o[18]~57 ;
wire \u0_m0_wo0_mtree_add1_4_o[20]~58_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[20]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[9]~29 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[10]~31 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[11]~33 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[12]~34_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[11]~32_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[10]~30_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_0_o[10]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[9]~28 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[10]~30 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[11]~32 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[12]~34 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[13]~36 ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[14]~37_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[14]~q ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[8]~28 ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[9]~30 ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[10]~32 ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[11]~34 ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[12]~36 ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[13]~37_combout ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[13]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[13]~35_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[13]~q ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[12]~35_combout ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[12]~33_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[11]~33_combout ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[11]~31_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[10]~31_combout ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[10]~q ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[10]~29_combout ;
wire \u0_m0_wo0_mtree_mult1_20_sub_2_o[10]~q ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[9]~29_combout ;
wire \u0_m0_wo0_mtree_mult1_21_add_1_o[9]~q ;
wire \u0_m0_wo0_mtree_add0_10_o[9]~32 ;
wire \u0_m0_wo0_mtree_add0_10_o[10]~34 ;
wire \u0_m0_wo0_mtree_add0_10_o[11]~36 ;
wire \u0_m0_wo0_mtree_add0_10_o[12]~38 ;
wire \u0_m0_wo0_mtree_add0_10_o[13]~40 ;
wire \u0_m0_wo0_mtree_add0_10_o[14]~42 ;
wire \u0_m0_wo0_mtree_add0_10_o[15]~43_combout ;
wire \u0_m0_wo0_mtree_add0_10_o[15]~q ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[9]~28 ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[10]~30 ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[11]~32 ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[12]~34 ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[13]~36 ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[14]~37_combout ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[14]~q ;
wire \u0_m0_wo0_mtree_add0_10_o[14]~41_combout ;
wire \u0_m0_wo0_mtree_add0_10_o[14]~q ;
wire \u0_m0_wo0_mtree_add0_10_o[13]~39_combout ;
wire \u0_m0_wo0_mtree_add0_10_o[13]~q ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[13]~35_combout ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[13]~q ;
wire \u0_m0_wo0_mtree_add0_10_o[12]~37_combout ;
wire \u0_m0_wo0_mtree_add0_10_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[12]~33_combout ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[12]~q ;
wire \u0_m0_wo0_mtree_add0_10_o[11]~35_combout ;
wire \u0_m0_wo0_mtree_add0_10_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[11]~31_combout ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[11]~q ;
wire \u0_m0_wo0_mtree_add0_10_o[10]~33_combout ;
wire \u0_m0_wo0_mtree_add0_10_o[10]~q ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[10]~29_combout ;
wire \u0_m0_wo0_mtree_mult1_22_sub_1_o[10]~q ;
wire \u0_m0_wo0_mtree_add1_5_o[9]~36 ;
wire \u0_m0_wo0_mtree_add1_5_o[10]~38 ;
wire \u0_m0_wo0_mtree_add1_5_o[11]~40 ;
wire \u0_m0_wo0_mtree_add1_5_o[12]~42 ;
wire \u0_m0_wo0_mtree_add1_5_o[13]~44 ;
wire \u0_m0_wo0_mtree_add1_5_o[14]~46 ;
wire \u0_m0_wo0_mtree_add1_5_o[15]~48 ;
wire \u0_m0_wo0_mtree_add1_5_o[17]~49_combout ;
wire \u0_m0_wo0_mtree_add1_5_o[17]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[18]~56_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[18]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[17]~54_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[17]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[16]~52_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[16]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[15]~50_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[15]~q ;
wire \u0_m0_wo0_mtree_add1_5_o[15]~47_combout ;
wire \u0_m0_wo0_mtree_add1_5_o[15]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[14]~48_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[14]~q ;
wire \u0_m0_wo0_mtree_add1_5_o[14]~45_combout ;
wire \u0_m0_wo0_mtree_add1_5_o[14]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[13]~46_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[13]~q ;
wire \u0_m0_wo0_mtree_add1_5_o[13]~43_combout ;
wire \u0_m0_wo0_mtree_add1_5_o[13]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[12]~44_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[12]~q ;
wire \u0_m0_wo0_mtree_add1_5_o[12]~41_combout ;
wire \u0_m0_wo0_mtree_add1_5_o[12]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[11]~42_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[11]~q ;
wire \u0_m0_wo0_mtree_add1_5_o[11]~39_combout ;
wire \u0_m0_wo0_mtree_add1_5_o[11]~q ;
wire \u0_m0_wo0_mtree_add1_4_o[10]~40_combout ;
wire \u0_m0_wo0_mtree_add1_4_o[10]~q ;
wire \u0_m0_wo0_mtree_add1_5_o[10]~37_combout ;
wire \u0_m0_wo0_mtree_add1_5_o[10]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[9]~40 ;
wire \u0_m0_wo0_mtree_add2_2_o[10]~42 ;
wire \u0_m0_wo0_mtree_add2_2_o[11]~44 ;
wire \u0_m0_wo0_mtree_add2_2_o[12]~46 ;
wire \u0_m0_wo0_mtree_add2_2_o[13]~48 ;
wire \u0_m0_wo0_mtree_add2_2_o[14]~50 ;
wire \u0_m0_wo0_mtree_add2_2_o[15]~52 ;
wire \u0_m0_wo0_mtree_add2_2_o[16]~54 ;
wire \u0_m0_wo0_mtree_add2_2_o[17]~56 ;
wire \u0_m0_wo0_mtree_add2_2_o[18]~58 ;
wire \u0_m0_wo0_mtree_add2_2_o[19]~60 ;
wire \u0_m0_wo0_mtree_add2_2_o[20]~61_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[20]~q ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[9]~29 ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[10]~31 ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[11]~33 ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[12]~34_combout ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[12]~q ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[11]~32_combout ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[11]~q ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[10]~30_combout ;
wire \u0_m0_wo0_mtree_mult1_25_sub_0_o[10]~q ;
wire \u0_m0_wo0_mtree_add0_12_o[9]~33 ;
wire \u0_m0_wo0_mtree_add0_12_o[10]~35 ;
wire \u0_m0_wo0_mtree_add0_12_o[11]~37 ;
wire \u0_m0_wo0_mtree_add0_12_o[12]~39 ;
wire \u0_m0_wo0_mtree_add0_12_o[13]~40_combout ;
wire \u0_m0_wo0_mtree_add0_12_o[13]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[19]~59_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[19]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[18]~57_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[18]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[17]~55_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[17]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[16]~53_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[16]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[15]~51_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[15]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[14]~49_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[14]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[13]~47_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[13]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[12]~45_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[12]~q ;
wire \u0_m0_wo0_mtree_add0_12_o[12]~38_combout ;
wire \u0_m0_wo0_mtree_add0_12_o[12]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[11]~43_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[11]~q ;
wire \u0_m0_wo0_mtree_add0_12_o[11]~36_combout ;
wire \u0_m0_wo0_mtree_add0_12_o[11]~q ;
wire \u0_m0_wo0_mtree_add2_2_o[10]~41_combout ;
wire \u0_m0_wo0_mtree_add2_2_o[10]~q ;
wire \u0_m0_wo0_mtree_add0_12_o[10]~34_combout ;
wire \u0_m0_wo0_mtree_add0_12_o[10]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[9]~40 ;
wire \u0_m0_wo0_mtree_add3_1_o[10]~42 ;
wire \u0_m0_wo0_mtree_add3_1_o[11]~44 ;
wire \u0_m0_wo0_mtree_add3_1_o[12]~46 ;
wire \u0_m0_wo0_mtree_add3_1_o[13]~48 ;
wire \u0_m0_wo0_mtree_add3_1_o[14]~50 ;
wire \u0_m0_wo0_mtree_add3_1_o[15]~52 ;
wire \u0_m0_wo0_mtree_add3_1_o[16]~54 ;
wire \u0_m0_wo0_mtree_add3_1_o[17]~56 ;
wire \u0_m0_wo0_mtree_add3_1_o[18]~58 ;
wire \u0_m0_wo0_mtree_add3_1_o[19]~60 ;
wire \u0_m0_wo0_mtree_add3_1_o[20]~61_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[20]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[19]~59_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[19]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[19]~59_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[19]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[18]~57_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[18]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[18]~57_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[18]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[17]~55_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[17]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[17]~55_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[17]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[16]~53_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[16]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[16]~53_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[16]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[15]~51_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[15]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[15]~51_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[15]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[14]~49_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[14]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[14]~49_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[14]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[13]~47_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[13]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[13]~47_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[13]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[12]~45_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[12]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[12]~45_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[12]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[11]~43_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[11]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[11]~43_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[11]~q ;
wire \u0_m0_wo0_mtree_add3_0_o[10]~41_combout ;
wire \u0_m0_wo0_mtree_add3_0_o[10]~q ;
wire \u0_m0_wo0_mtree_add3_1_o[10]~41_combout ;
wire \u0_m0_wo0_mtree_add3_1_o[10]~q ;
wire \u0_m0_wo0_mtree_add4_0_o[9]~31 ;
wire \u0_m0_wo0_mtree_add4_0_o[10]~33 ;
wire \u0_m0_wo0_mtree_add4_0_o[11]~35 ;
wire \u0_m0_wo0_mtree_add4_0_o[12]~37 ;
wire \u0_m0_wo0_mtree_add4_0_o[13]~39 ;
wire \u0_m0_wo0_mtree_add4_0_o[14]~41 ;
wire \u0_m0_wo0_mtree_add4_0_o[15]~43 ;
wire \u0_m0_wo0_mtree_add4_0_o[16]~45 ;
wire \u0_m0_wo0_mtree_add4_0_o[17]~47 ;
wire \u0_m0_wo0_mtree_add4_0_o[18]~49 ;
wire \u0_m0_wo0_mtree_add4_0_o[19]~51 ;
wire \u0_m0_wo0_mtree_add4_0_o[20]~52_combout ;
wire \u0_m0_wo0_mtree_add4_0_o[19]~50_combout ;
wire \u0_m0_wo0_mtree_add4_0_o[18]~48_combout ;
wire \u0_m0_wo0_mtree_add4_0_o[17]~46_combout ;
wire \u0_m0_wo0_mtree_add4_0_o[16]~44_combout ;
wire \u0_m0_wo0_mtree_add4_0_o[15]~42_combout ;
wire \u0_m0_wo0_mtree_add4_0_o[14]~40_combout ;
wire \u0_m0_wo0_mtree_add4_0_o[13]~38_combout ;
wire \u0_m0_wo0_mtree_add4_0_o[12]~36_combout ;
wire \u0_m0_wo0_mtree_add4_0_o[11]~34_combout ;
wire \u0_m0_wo0_mtree_add4_0_o[10]~32_combout ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[9]~29 ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[10]~31 ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[11]~33 ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[12]~34_combout ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[11]~32_combout ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[10]~30_combout ;
wire \u1_m0_wo0_mtree_mult1_5_sub_0_o[10]~q ;
wire \u1_m0_wo0_mtree_add1_1_o[9]~33 ;
wire \u1_m0_wo0_mtree_add1_1_o[10]~35 ;
wire \u1_m0_wo0_mtree_add1_1_o[11]~37 ;
wire \u1_m0_wo0_mtree_add1_1_o[12]~39 ;
wire \u1_m0_wo0_mtree_add1_1_o[15]~40_combout ;
wire \u1_m0_wo0_mtree_add1_1_o[15]~q ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[9]~28 ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[10]~30 ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[11]~32 ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[12]~34 ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[13]~36 ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[14]~37_combout ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[14]~q ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[8]~28 ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[9]~30 ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[10]~32 ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[11]~34 ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[12]~36 ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[13]~37_combout ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[13]~q ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[13]~35_combout ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[13]~q ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[12]~35_combout ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[12]~33_combout ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[11]~33_combout ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[11]~31_combout ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[10]~31_combout ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[10]~q ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[10]~29_combout ;
wire \u1_m0_wo0_mtree_mult1_8_sub_1_o[10]~q ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[9]~29_combout ;
wire \u1_m0_wo0_mtree_mult1_9_add_1_o[9]~q ;
wire \u1_m0_wo0_mtree_add0_4_o[9]~32 ;
wire \u1_m0_wo0_mtree_add0_4_o[10]~34 ;
wire \u1_m0_wo0_mtree_add0_4_o[11]~36 ;
wire \u1_m0_wo0_mtree_add0_4_o[12]~38 ;
wire \u1_m0_wo0_mtree_add0_4_o[13]~40 ;
wire \u1_m0_wo0_mtree_add0_4_o[14]~42 ;
wire \u1_m0_wo0_mtree_add0_4_o[15]~43_combout ;
wire \u1_m0_wo0_mtree_add0_4_o[15]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[9]~29 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[10]~31 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[11]~33 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[12]~34_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[11]~32_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[10]~30_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_0_o[10]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[9]~28 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[10]~30 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[11]~32 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[12]~34 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[13]~36 ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[14]~37_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[14]~q ;
wire \u1_m0_wo0_mtree_add0_4_o[14]~41_combout ;
wire \u1_m0_wo0_mtree_add0_4_o[14]~q ;
wire \u1_m0_wo0_mtree_add0_4_o[13]~39_combout ;
wire \u1_m0_wo0_mtree_add0_4_o[13]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[13]~35_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[13]~q ;
wire \u1_m0_wo0_mtree_add0_4_o[12]~37_combout ;
wire \u1_m0_wo0_mtree_add0_4_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[12]~33_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[12]~q ;
wire \u1_m0_wo0_mtree_add0_4_o[11]~35_combout ;
wire \u1_m0_wo0_mtree_add0_4_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[11]~31_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[11]~q ;
wire \u1_m0_wo0_mtree_add0_4_o[10]~33_combout ;
wire \u1_m0_wo0_mtree_add0_4_o[10]~q ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[10]~29_combout ;
wire \u1_m0_wo0_mtree_mult1_10_sub_2_o[10]~q ;
wire \u1_m0_wo0_mtree_add1_2_o[9]~36 ;
wire \u1_m0_wo0_mtree_add1_2_o[10]~38 ;
wire \u1_m0_wo0_mtree_add1_2_o[11]~40 ;
wire \u1_m0_wo0_mtree_add1_2_o[12]~42 ;
wire \u1_m0_wo0_mtree_add1_2_o[13]~44 ;
wire \u1_m0_wo0_mtree_add1_2_o[14]~46 ;
wire \u1_m0_wo0_mtree_add1_2_o[15]~48 ;
wire \u1_m0_wo0_mtree_add1_2_o[17]~49_combout ;
wire \u1_m0_wo0_mtree_add1_2_o[17]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[9]~30 ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[10]~32 ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[11]~34 ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[12]~36 ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[13]~37_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[13]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[12]~35_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[11]~33_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[10]~31_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_1_o[10]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[9]~26 ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[10]~28 ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[11]~30 ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[12]~32 ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[13]~34 ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[14]~36 ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[15]~37_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[15]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[9]~32 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[10]~34 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[11]~36 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[12]~38 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[13]~40 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[14]~42 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[15]~43_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[15]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[14]~41_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[14]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[13]~39_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[13]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[12]~37_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[11]~35_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[10]~33_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_1_o[10]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[9]~22 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[10]~24 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[11]~26 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[12]~28 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[13]~30 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[14]~32 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[15]~34 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[16]~36 ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[17]~37_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[17]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[16]~35_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[16]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[15]~33_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[15]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[14]~35_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[14]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[14]~31_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[14]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[13]~33_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[13]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[13]~29_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[13]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[12]~31_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[12]~27_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[11]~29_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[11]~25_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[10]~27_combout ;
wire \u1_m0_wo0_mtree_mult1_12_add_3_o[10]~q ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[10]~23_combout ;
wire \u1_m0_wo0_mtree_mult1_13_sub_3_o[10]~q ;
wire \u1_m0_wo0_mtree_add0_6_o[9]~38 ;
wire \u1_m0_wo0_mtree_add0_6_o[10]~40 ;
wire \u1_m0_wo0_mtree_add0_6_o[11]~42 ;
wire \u1_m0_wo0_mtree_add0_6_o[12]~44 ;
wire \u1_m0_wo0_mtree_add0_6_o[13]~46 ;
wire \u1_m0_wo0_mtree_add0_6_o[14]~48 ;
wire \u1_m0_wo0_mtree_add0_6_o[15]~50 ;
wire \u1_m0_wo0_mtree_add0_6_o[16]~52 ;
wire \u1_m0_wo0_mtree_add0_6_o[17]~54 ;
wire \u1_m0_wo0_mtree_add0_6_o[18]~55_combout ;
wire \u1_m0_wo0_mtree_add0_6_o[18]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[9]~28 ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[10]~30 ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[11]~32 ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[12]~34 ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[13]~36 ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[14]~37_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[14]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[13]~35_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[13]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[12]~33_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[11]~31_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[10]~29_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_1_o[10]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[9]~22 ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[10]~24 ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[11]~26 ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[12]~28 ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[13]~30 ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[14]~32 ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[15]~34 ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[16]~36 ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[17]~37_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[17]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[9]~36 ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[10]~38 ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[11]~40 ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[12]~42 ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[13]~44 ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[14]~46 ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[15]~48 ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[16]~50 ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[17]~52 ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[18]~54 ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[19]~55_combout ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[19]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[18]~53_combout ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[18]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[17]~51_combout ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[17]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[16]~35_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[16]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[16]~49_combout ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[16]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[15]~33_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[15]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[15]~47_combout ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[15]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[14]~31_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[14]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[14]~45_combout ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[14]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[13]~29_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[13]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[13]~43_combout ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[13]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[12]~27_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[12]~41_combout ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[11]~25_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[11]~39_combout ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[10]~23_combout ;
wire \u1_m0_wo0_mtree_mult1_14_add_3_o[10]~q ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[10]~37_combout ;
wire \u1_m0_wo0_mtree_mult1_15_sub_1_o[10]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[9]~40 ;
wire \u1_m0_wo0_mtree_add0_7_o[10]~42 ;
wire \u1_m0_wo0_mtree_add0_7_o[11]~44 ;
wire \u1_m0_wo0_mtree_add0_7_o[12]~46 ;
wire \u1_m0_wo0_mtree_add0_7_o[13]~48 ;
wire \u1_m0_wo0_mtree_add0_7_o[14]~50 ;
wire \u1_m0_wo0_mtree_add0_7_o[15]~52 ;
wire \u1_m0_wo0_mtree_add0_7_o[16]~54 ;
wire \u1_m0_wo0_mtree_add0_7_o[17]~56 ;
wire \u1_m0_wo0_mtree_add0_7_o[18]~58 ;
wire \u1_m0_wo0_mtree_add0_7_o[19]~60 ;
wire \u1_m0_wo0_mtree_add0_7_o[20]~61_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[20]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[19]~59_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[19]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[18]~57_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[18]~q ;
wire \u1_m0_wo0_mtree_add0_6_o[17]~53_combout ;
wire \u1_m0_wo0_mtree_add0_6_o[17]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[17]~55_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[17]~q ;
wire \u1_m0_wo0_mtree_add0_6_o[16]~51_combout ;
wire \u1_m0_wo0_mtree_add0_6_o[16]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[16]~53_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[16]~q ;
wire \u1_m0_wo0_mtree_add0_6_o[15]~49_combout ;
wire \u1_m0_wo0_mtree_add0_6_o[15]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[15]~51_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[15]~q ;
wire \u1_m0_wo0_mtree_add0_6_o[14]~47_combout ;
wire \u1_m0_wo0_mtree_add0_6_o[14]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[14]~49_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[14]~q ;
wire \u1_m0_wo0_mtree_add0_6_o[13]~45_combout ;
wire \u1_m0_wo0_mtree_add0_6_o[13]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[13]~47_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[13]~q ;
wire \u1_m0_wo0_mtree_add0_6_o[12]~43_combout ;
wire \u1_m0_wo0_mtree_add0_6_o[12]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[12]~45_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[12]~q ;
wire \u1_m0_wo0_mtree_add0_6_o[11]~41_combout ;
wire \u1_m0_wo0_mtree_add0_6_o[11]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[11]~43_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[11]~q ;
wire \u1_m0_wo0_mtree_add0_6_o[10]~39_combout ;
wire \u1_m0_wo0_mtree_add0_6_o[10]~q ;
wire \u1_m0_wo0_mtree_add0_7_o[10]~41_combout ;
wire \u1_m0_wo0_mtree_add0_7_o[10]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[9]~40 ;
wire \u1_m0_wo0_mtree_add1_3_o[10]~42 ;
wire \u1_m0_wo0_mtree_add1_3_o[11]~44 ;
wire \u1_m0_wo0_mtree_add1_3_o[12]~46 ;
wire \u1_m0_wo0_mtree_add1_3_o[13]~48 ;
wire \u1_m0_wo0_mtree_add1_3_o[14]~50 ;
wire \u1_m0_wo0_mtree_add1_3_o[15]~52 ;
wire \u1_m0_wo0_mtree_add1_3_o[16]~54 ;
wire \u1_m0_wo0_mtree_add1_3_o[17]~56 ;
wire \u1_m0_wo0_mtree_add1_3_o[18]~58 ;
wire \u1_m0_wo0_mtree_add1_3_o[19]~60 ;
wire \u1_m0_wo0_mtree_add1_3_o[20]~61_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[20]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[19]~59_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[19]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[18]~57_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[18]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[17]~55_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[17]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[16]~53_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[16]~q ;
wire \u1_m0_wo0_mtree_add1_2_o[15]~47_combout ;
wire \u1_m0_wo0_mtree_add1_2_o[15]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[15]~51_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[15]~q ;
wire \u1_m0_wo0_mtree_add1_2_o[14]~45_combout ;
wire \u1_m0_wo0_mtree_add1_2_o[14]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[14]~49_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[14]~q ;
wire \u1_m0_wo0_mtree_add1_2_o[13]~43_combout ;
wire \u1_m0_wo0_mtree_add1_2_o[13]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[13]~47_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[13]~q ;
wire \u1_m0_wo0_mtree_add1_2_o[12]~41_combout ;
wire \u1_m0_wo0_mtree_add1_2_o[12]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[12]~45_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[12]~q ;
wire \u1_m0_wo0_mtree_add1_2_o[11]~39_combout ;
wire \u1_m0_wo0_mtree_add1_2_o[11]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[11]~43_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[11]~q ;
wire \u1_m0_wo0_mtree_add1_2_o[10]~37_combout ;
wire \u1_m0_wo0_mtree_add1_2_o[10]~q ;
wire \u1_m0_wo0_mtree_add1_3_o[10]~41_combout ;
wire \u1_m0_wo0_mtree_add1_3_o[10]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[9]~40 ;
wire \u1_m0_wo0_mtree_add2_1_o[10]~42 ;
wire \u1_m0_wo0_mtree_add2_1_o[11]~44 ;
wire \u1_m0_wo0_mtree_add2_1_o[12]~46 ;
wire \u1_m0_wo0_mtree_add2_1_o[13]~48 ;
wire \u1_m0_wo0_mtree_add2_1_o[14]~50 ;
wire \u1_m0_wo0_mtree_add2_1_o[15]~52 ;
wire \u1_m0_wo0_mtree_add2_1_o[16]~54 ;
wire \u1_m0_wo0_mtree_add2_1_o[17]~56 ;
wire \u1_m0_wo0_mtree_add2_1_o[18]~58 ;
wire \u1_m0_wo0_mtree_add2_1_o[19]~60 ;
wire \u1_m0_wo0_mtree_add2_1_o[20]~61_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[20]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[19]~59_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[19]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[18]~57_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[18]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[17]~55_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[17]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[16]~53_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[16]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[15]~51_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[15]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[14]~49_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[14]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[13]~47_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[13]~q ;
wire \u1_m0_wo0_mtree_add1_1_o[12]~38_combout ;
wire \u1_m0_wo0_mtree_add1_1_o[12]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[12]~45_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[12]~q ;
wire \u1_m0_wo0_mtree_add1_1_o[11]~36_combout ;
wire \u1_m0_wo0_mtree_add1_1_o[11]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[11]~43_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[11]~q ;
wire \u1_m0_wo0_mtree_add1_1_o[10]~34_combout ;
wire \u1_m0_wo0_mtree_add1_1_o[10]~q ;
wire \u1_m0_wo0_mtree_add2_1_o[10]~41_combout ;
wire \u1_m0_wo0_mtree_add2_1_o[10]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[9]~40 ;
wire \u1_m0_wo0_mtree_add3_0_o[10]~42 ;
wire \u1_m0_wo0_mtree_add3_0_o[11]~44 ;
wire \u1_m0_wo0_mtree_add3_0_o[12]~46 ;
wire \u1_m0_wo0_mtree_add3_0_o[13]~48 ;
wire \u1_m0_wo0_mtree_add3_0_o[14]~50 ;
wire \u1_m0_wo0_mtree_add3_0_o[15]~52 ;
wire \u1_m0_wo0_mtree_add3_0_o[16]~54 ;
wire \u1_m0_wo0_mtree_add3_0_o[17]~56 ;
wire \u1_m0_wo0_mtree_add3_0_o[18]~58 ;
wire \u1_m0_wo0_mtree_add3_0_o[19]~60 ;
wire \u1_m0_wo0_mtree_add3_0_o[20]~61_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[20]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[9]~28 ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[10]~30 ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[11]~32 ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[12]~34 ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[13]~36 ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[14]~37_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[14]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[13]~35_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[13]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[12]~33_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[11]~31_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[10]~29_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_1_o[10]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[9]~22 ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[10]~24 ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[11]~26 ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[12]~28 ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[13]~30 ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[14]~32 ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[15]~34 ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[16]~36 ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[17]~37_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[17]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[9]~32 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[10]~34 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[11]~36 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[12]~38 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[13]~40 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[14]~42 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[15]~43_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[15]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[14]~41_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[14]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[13]~39_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[13]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[12]~37_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[11]~35_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[10]~33_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_1_o[10]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[9]~22 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[10]~24 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[11]~26 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[12]~28 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[13]~30 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[14]~32 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[15]~34 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[16]~36 ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[17]~37_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[17]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[16]~35_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[16]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[16]~35_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[16]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[15]~33_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[15]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[15]~33_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[15]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[14]~31_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[14]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[14]~31_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[14]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[13]~29_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[13]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[13]~29_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[13]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[12]~27_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[12]~27_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[11]~25_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[11]~25_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[10]~23_combout ;
wire \u1_m0_wo0_mtree_mult1_16_add_3_o[10]~q ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[10]~23_combout ;
wire \u1_m0_wo0_mtree_mult1_17_sub_3_o[10]~q ;
wire \u1_m0_wo0_mtree_add0_8_o[9]~38 ;
wire \u1_m0_wo0_mtree_add0_8_o[10]~40 ;
wire \u1_m0_wo0_mtree_add0_8_o[11]~42 ;
wire \u1_m0_wo0_mtree_add0_8_o[12]~44 ;
wire \u1_m0_wo0_mtree_add0_8_o[13]~46 ;
wire \u1_m0_wo0_mtree_add0_8_o[14]~48 ;
wire \u1_m0_wo0_mtree_add0_8_o[15]~50 ;
wire \u1_m0_wo0_mtree_add0_8_o[16]~52 ;
wire \u1_m0_wo0_mtree_add0_8_o[17]~54 ;
wire \u1_m0_wo0_mtree_add0_8_o[18]~55_combout ;
wire \u1_m0_wo0_mtree_add0_8_o[18]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[9]~30 ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[10]~32 ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[11]~34 ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[12]~36 ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[13]~37_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[13]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[12]~35_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[11]~33_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[10]~31_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_1_o[10]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[9]~26 ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[10]~28 ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[11]~30 ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[12]~32 ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[13]~34 ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[14]~36 ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[15]~37_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[15]~q ;
wire \u1_m0_wo0_mtree_add0_8_o[17]~53_combout ;
wire \u1_m0_wo0_mtree_add0_8_o[17]~q ;
wire \u1_m0_wo0_mtree_add0_8_o[16]~51_combout ;
wire \u1_m0_wo0_mtree_add0_8_o[16]~q ;
wire \u1_m0_wo0_mtree_add0_8_o[15]~49_combout ;
wire \u1_m0_wo0_mtree_add0_8_o[15]~q ;
wire \u1_m0_wo0_mtree_add0_8_o[14]~47_combout ;
wire \u1_m0_wo0_mtree_add0_8_o[14]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[14]~35_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[14]~q ;
wire \u1_m0_wo0_mtree_add0_8_o[13]~45_combout ;
wire \u1_m0_wo0_mtree_add0_8_o[13]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[13]~33_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[13]~q ;
wire \u1_m0_wo0_mtree_add0_8_o[12]~43_combout ;
wire \u1_m0_wo0_mtree_add0_8_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[12]~31_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[12]~q ;
wire \u1_m0_wo0_mtree_add0_8_o[11]~41_combout ;
wire \u1_m0_wo0_mtree_add0_8_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[11]~29_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[11]~q ;
wire \u1_m0_wo0_mtree_add0_8_o[10]~39_combout ;
wire \u1_m0_wo0_mtree_add0_8_o[10]~q ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[10]~27_combout ;
wire \u1_m0_wo0_mtree_mult1_18_add_3_o[10]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[9]~39 ;
wire \u1_m0_wo0_mtree_add1_4_o[10]~41 ;
wire \u1_m0_wo0_mtree_add1_4_o[11]~43 ;
wire \u1_m0_wo0_mtree_add1_4_o[12]~45 ;
wire \u1_m0_wo0_mtree_add1_4_o[13]~47 ;
wire \u1_m0_wo0_mtree_add1_4_o[14]~49 ;
wire \u1_m0_wo0_mtree_add1_4_o[15]~51 ;
wire \u1_m0_wo0_mtree_add1_4_o[16]~53 ;
wire \u1_m0_wo0_mtree_add1_4_o[17]~55 ;
wire \u1_m0_wo0_mtree_add1_4_o[18]~57 ;
wire \u1_m0_wo0_mtree_add1_4_o[20]~58_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[20]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[9]~29 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[10]~31 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[11]~33 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[12]~34_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[11]~32_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[10]~30_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_0_o[10]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[9]~28 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[10]~30 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[11]~32 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[12]~34 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[13]~36 ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[14]~37_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[14]~q ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[8]~28 ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[9]~30 ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[10]~32 ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[11]~34 ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[12]~36 ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[13]~37_combout ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[13]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[13]~35_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[13]~q ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[12]~35_combout ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[12]~33_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[11]~33_combout ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[11]~31_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[10]~31_combout ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[10]~q ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[10]~29_combout ;
wire \u1_m0_wo0_mtree_mult1_20_sub_2_o[10]~q ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[9]~29_combout ;
wire \u1_m0_wo0_mtree_mult1_21_add_1_o[9]~q ;
wire \u1_m0_wo0_mtree_add0_10_o[9]~32 ;
wire \u1_m0_wo0_mtree_add0_10_o[10]~34 ;
wire \u1_m0_wo0_mtree_add0_10_o[11]~36 ;
wire \u1_m0_wo0_mtree_add0_10_o[12]~38 ;
wire \u1_m0_wo0_mtree_add0_10_o[13]~40 ;
wire \u1_m0_wo0_mtree_add0_10_o[14]~42 ;
wire \u1_m0_wo0_mtree_add0_10_o[15]~43_combout ;
wire \u1_m0_wo0_mtree_add0_10_o[15]~q ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[9]~28 ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[10]~30 ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[11]~32 ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[12]~34 ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[13]~36 ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[14]~37_combout ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[14]~q ;
wire \u1_m0_wo0_mtree_add0_10_o[14]~41_combout ;
wire \u1_m0_wo0_mtree_add0_10_o[14]~q ;
wire \u1_m0_wo0_mtree_add0_10_o[13]~39_combout ;
wire \u1_m0_wo0_mtree_add0_10_o[13]~q ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[13]~35_combout ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[13]~q ;
wire \u1_m0_wo0_mtree_add0_10_o[12]~37_combout ;
wire \u1_m0_wo0_mtree_add0_10_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[12]~33_combout ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[12]~q ;
wire \u1_m0_wo0_mtree_add0_10_o[11]~35_combout ;
wire \u1_m0_wo0_mtree_add0_10_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[11]~31_combout ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[11]~q ;
wire \u1_m0_wo0_mtree_add0_10_o[10]~33_combout ;
wire \u1_m0_wo0_mtree_add0_10_o[10]~q ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[10]~29_combout ;
wire \u1_m0_wo0_mtree_mult1_22_sub_1_o[10]~q ;
wire \u1_m0_wo0_mtree_add1_5_o[9]~36 ;
wire \u1_m0_wo0_mtree_add1_5_o[10]~38 ;
wire \u1_m0_wo0_mtree_add1_5_o[11]~40 ;
wire \u1_m0_wo0_mtree_add1_5_o[12]~42 ;
wire \u1_m0_wo0_mtree_add1_5_o[13]~44 ;
wire \u1_m0_wo0_mtree_add1_5_o[14]~46 ;
wire \u1_m0_wo0_mtree_add1_5_o[15]~48 ;
wire \u1_m0_wo0_mtree_add1_5_o[17]~49_combout ;
wire \u1_m0_wo0_mtree_add1_5_o[17]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[18]~56_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[18]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[17]~54_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[17]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[16]~52_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[16]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[15]~50_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[15]~q ;
wire \u1_m0_wo0_mtree_add1_5_o[15]~47_combout ;
wire \u1_m0_wo0_mtree_add1_5_o[15]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[14]~48_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[14]~q ;
wire \u1_m0_wo0_mtree_add1_5_o[14]~45_combout ;
wire \u1_m0_wo0_mtree_add1_5_o[14]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[13]~46_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[13]~q ;
wire \u1_m0_wo0_mtree_add1_5_o[13]~43_combout ;
wire \u1_m0_wo0_mtree_add1_5_o[13]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[12]~44_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[12]~q ;
wire \u1_m0_wo0_mtree_add1_5_o[12]~41_combout ;
wire \u1_m0_wo0_mtree_add1_5_o[12]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[11]~42_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[11]~q ;
wire \u1_m0_wo0_mtree_add1_5_o[11]~39_combout ;
wire \u1_m0_wo0_mtree_add1_5_o[11]~q ;
wire \u1_m0_wo0_mtree_add1_4_o[10]~40_combout ;
wire \u1_m0_wo0_mtree_add1_4_o[10]~q ;
wire \u1_m0_wo0_mtree_add1_5_o[10]~37_combout ;
wire \u1_m0_wo0_mtree_add1_5_o[10]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[9]~40 ;
wire \u1_m0_wo0_mtree_add2_2_o[10]~42 ;
wire \u1_m0_wo0_mtree_add2_2_o[11]~44 ;
wire \u1_m0_wo0_mtree_add2_2_o[12]~46 ;
wire \u1_m0_wo0_mtree_add2_2_o[13]~48 ;
wire \u1_m0_wo0_mtree_add2_2_o[14]~50 ;
wire \u1_m0_wo0_mtree_add2_2_o[15]~52 ;
wire \u1_m0_wo0_mtree_add2_2_o[16]~54 ;
wire \u1_m0_wo0_mtree_add2_2_o[17]~56 ;
wire \u1_m0_wo0_mtree_add2_2_o[18]~58 ;
wire \u1_m0_wo0_mtree_add2_2_o[19]~60 ;
wire \u1_m0_wo0_mtree_add2_2_o[20]~61_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[20]~q ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[9]~29 ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[10]~31 ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[11]~33 ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[12]~34_combout ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[12]~q ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[11]~32_combout ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[11]~q ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[10]~30_combout ;
wire \u1_m0_wo0_mtree_mult1_25_sub_0_o[10]~q ;
wire \u1_m0_wo0_mtree_add0_12_o[9]~33 ;
wire \u1_m0_wo0_mtree_add0_12_o[10]~35 ;
wire \u1_m0_wo0_mtree_add0_12_o[11]~37 ;
wire \u1_m0_wo0_mtree_add0_12_o[12]~39 ;
wire \u1_m0_wo0_mtree_add0_12_o[13]~40_combout ;
wire \u1_m0_wo0_mtree_add0_12_o[13]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[19]~59_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[19]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[18]~57_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[18]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[17]~55_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[17]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[16]~53_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[16]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[15]~51_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[15]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[14]~49_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[14]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[13]~47_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[13]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[12]~45_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[12]~q ;
wire \u1_m0_wo0_mtree_add0_12_o[12]~38_combout ;
wire \u1_m0_wo0_mtree_add0_12_o[12]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[11]~43_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[11]~q ;
wire \u1_m0_wo0_mtree_add0_12_o[11]~36_combout ;
wire \u1_m0_wo0_mtree_add0_12_o[11]~q ;
wire \u1_m0_wo0_mtree_add2_2_o[10]~41_combout ;
wire \u1_m0_wo0_mtree_add2_2_o[10]~q ;
wire \u1_m0_wo0_mtree_add0_12_o[10]~34_combout ;
wire \u1_m0_wo0_mtree_add0_12_o[10]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[9]~40 ;
wire \u1_m0_wo0_mtree_add3_1_o[10]~42 ;
wire \u1_m0_wo0_mtree_add3_1_o[11]~44 ;
wire \u1_m0_wo0_mtree_add3_1_o[12]~46 ;
wire \u1_m0_wo0_mtree_add3_1_o[13]~48 ;
wire \u1_m0_wo0_mtree_add3_1_o[14]~50 ;
wire \u1_m0_wo0_mtree_add3_1_o[15]~52 ;
wire \u1_m0_wo0_mtree_add3_1_o[16]~54 ;
wire \u1_m0_wo0_mtree_add3_1_o[17]~56 ;
wire \u1_m0_wo0_mtree_add3_1_o[18]~58 ;
wire \u1_m0_wo0_mtree_add3_1_o[19]~60 ;
wire \u1_m0_wo0_mtree_add3_1_o[20]~61_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[20]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[19]~59_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[19]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[19]~59_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[19]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[18]~57_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[18]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[18]~57_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[18]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[17]~55_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[17]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[17]~55_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[17]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[16]~53_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[16]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[16]~53_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[16]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[15]~51_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[15]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[15]~51_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[15]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[14]~49_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[14]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[14]~49_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[14]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[13]~47_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[13]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[13]~47_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[13]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[12]~45_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[12]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[12]~45_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[12]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[11]~43_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[11]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[11]~43_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[11]~q ;
wire \u1_m0_wo0_mtree_add3_0_o[10]~41_combout ;
wire \u1_m0_wo0_mtree_add3_0_o[10]~q ;
wire \u1_m0_wo0_mtree_add3_1_o[10]~41_combout ;
wire \u1_m0_wo0_mtree_add3_1_o[10]~q ;
wire \u1_m0_wo0_mtree_add4_0_o[9]~31 ;
wire \u1_m0_wo0_mtree_add4_0_o[10]~33 ;
wire \u1_m0_wo0_mtree_add4_0_o[11]~35 ;
wire \u1_m0_wo0_mtree_add4_0_o[12]~37 ;
wire \u1_m0_wo0_mtree_add4_0_o[13]~39 ;
wire \u1_m0_wo0_mtree_add4_0_o[14]~41 ;
wire \u1_m0_wo0_mtree_add4_0_o[15]~43 ;
wire \u1_m0_wo0_mtree_add4_0_o[16]~45 ;
wire \u1_m0_wo0_mtree_add4_0_o[17]~47 ;
wire \u1_m0_wo0_mtree_add4_0_o[18]~49 ;
wire \u1_m0_wo0_mtree_add4_0_o[19]~51 ;
wire \u1_m0_wo0_mtree_add4_0_o[20]~52_combout ;
wire \u1_m0_wo0_mtree_add4_0_o[19]~50_combout ;
wire \u1_m0_wo0_mtree_add4_0_o[18]~48_combout ;
wire \u1_m0_wo0_mtree_add4_0_o[17]~46_combout ;
wire \u1_m0_wo0_mtree_add4_0_o[16]~44_combout ;
wire \u1_m0_wo0_mtree_add4_0_o[15]~42_combout ;
wire \u1_m0_wo0_mtree_add4_0_o[14]~40_combout ;
wire \u1_m0_wo0_mtree_add4_0_o[13]~38_combout ;
wire \u1_m0_wo0_mtree_add4_0_o[12]~36_combout ;
wire \u1_m0_wo0_mtree_add4_0_o[11]~34_combout ;
wire \u1_m0_wo0_mtree_add4_0_o[10]~32_combout ;


lms_dsp_dspba_delay_2 d_u0_m0_wo0_compute_q_16(
	.aclr(areset),
	.delay_signals_0_0(\d_u0_m0_wo0_compute_q_16|delay_signals[0][0]~q ),
	.xin({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\d_u0_m0_wo0_compute_q_13|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_54 u0_m0_wo0_wi0_r0_delayr25(
	.aclr(areset),
	.xin({\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][0]~q }),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][2]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][0]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][1]~q ),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][10]~q ),
	.ena(\d_u0_m0_wo0_compute_q_13|delay_signals[0][0]~q ),
	.clk(clk));

lms_dsp_dspba_delay_16 d_u0_m0_wo0_wi0_r0_delayr24_q_14(
	.aclr(areset),
	.delay_signals_9_0(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][1]~q ),
	.delay_signals_0_0(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][0]~q ),
	.delay_signals_11_0(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][10]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_53 u0_m0_wo0_wi0_r0_delayr24(
	.aclr(areset),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][0]~q ),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr24|delay_signals[0][10]~q ),
	.ena(\d_u0_m0_wo0_compute_q_13|delay_signals[0][0]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_52 u0_m0_wo0_wi0_r0_delayr23(
	.aclr(areset),
	.xin({\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][11]~q ,\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][10]~q ,\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][9]~q ,\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][8]~q ,
\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][7]~q ,\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][6]~q ,\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][5]~q ,\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][4]~q ,
\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][3]~q ,\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][2]~q ,\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][1]~q ,\u0_m0_wo0_mtree_add0_4_o[0]~q }),
	.ena(\d_u0_m0_wo0_compute_q_13|delay_signals[0][0]~q ),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][0]~q ),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr23|delay_signals[0][10]~q ),
	.clk(clk));

lms_dsp_dspba_delay_15 d_u0_m0_wo0_wi0_r0_delayr22_q_13(
	.aclr(areset),
	.u0_m0_wo0_mtree_mult1_8_sub_1_o_1(\u0_m0_wo0_mtree_mult1_8_sub_1_o[1]~q ),
	.delay_signals_9_0(\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][1]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][2]~q ,gnd,gnd}),
	.delay_signals_11_0(\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u0_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][10]~q ),
	.clk(clk));

lms_dsp_dspba_delay_51 u0_m0_wo0_wi0_r0_delayr22(
	.aclr(areset),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][7]~q ),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][9]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][6]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][8]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][0]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][0]~q }),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][10]~q ),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][11]~q ),
	.ena(\d_u0_m0_wo0_compute_q_11|delay_signals[0][0]~q ),
	.clk(clk));

lms_dsp_dspba_delay_50 u0_m0_wo0_wi0_r0_delayr21(
	.aclr(areset),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][0]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][0]~q }),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][10]~q ),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][9]~q ),
	.ena(\d_u0_m0_wo0_compute_q_11|delay_signals[0][0]~q ),
	.clk(clk));

lms_dsp_dspba_delay_14 d_u0_m0_wo0_wi0_r0_delayr20_q_12(
	.aclr(areset),
	.delay_signals_7_0(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][1]~q ),
	.delay_signals_11_0(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][10]~q ),
	.delay_signals_9_0(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][8]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][1]~q ,gnd}),
	.clk(clk));

lms_dsp_dspba_delay_49 u0_m0_wo0_wi0_r0_delayr20(
	.aclr(areset),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][7]~q ),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][8]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][2]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][0]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][1]~q ),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][10]~q ),
	.ena(\d_u0_m0_wo0_compute_q_11|delay_signals[0][0]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_47 u0_m0_wo0_wi0_r0_delayr19(
	.aclr(areset),
	.xin({\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][11]~q ,\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][10]~q ,\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][9]~q ,\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][8]~q ,
\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][7]~q ,\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][6]~q ,\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][5]~q ,\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][4]~q ,
\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][3]~q ,\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][2]~q ,\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][1]~q ,\u0_m0_wo0_mtree_mult1_12_add_1_o[0]~q }),
	.ena(\d_u0_m0_wo0_compute_q_11|delay_signals[0][0]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][7]~q ),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][8]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][2]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][0]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][1]~q ),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr19|delay_signals[0][10]~q ),
	.clk(clk));

lms_dsp_dspba_delay_13 d_u0_m0_wo0_wi0_r0_delayr18_q_11(
	.aclr(areset),
	.delay_signals_6_0(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][1]~q ),
	.delay_signals_11_0(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][10]~q ),
	.delay_signals_9_0(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][7]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][1]~q ,gnd}),
	.clk(clk));

lms_dsp_dspba_delay_46 u0_m0_wo0_wi0_r0_delayr18(
	.aclr(areset),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][6]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][8]~q ),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][9]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][7]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][0]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][0]~q }),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][10]~q ),
	.ena(xIn_v[0]),
	.clk(clk));

lms_dsp_dspba_delay_12 d_u0_m0_wo0_wi0_r0_delayr17_q_11(
	.aclr(areset),
	.delay_signals_4_0(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][1]~q ),
	.delay_signals_11_0(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][10]~q ),
	.delay_signals_9_0(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][5]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][1]~q ,gnd}),
	.clk(clk));

lms_dsp_dspba_delay_45 u0_m0_wo0_wi0_r0_delayr17(
	.aclr(areset),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][4]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][6]~q ),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][9]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][5]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][7]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][0]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][0]~q }),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][10]~q ),
	.ena(xIn_v[0]),
	.clk(clk));

lms_dsp_dspba_delay_11 d_u0_m0_wo0_wi0_r0_delayr16_q_11(
	.aclr(areset),
	.delay_signals_4_0(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][2]~q ),
	.delay_signals_11_0(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][10]~q ),
	.delay_signals_9_0(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][5]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][2]~q ,gnd,gnd}),
	.clk(clk));

lms_dsp_dspba_delay_44 u0_m0_wo0_wi0_r0_delayr16(
	.aclr(areset),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][4]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][7]~q ),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][9]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][6]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][8]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][5]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][0]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][0]~q }),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][10]~q ),
	.ena(xIn_v[0]),
	.clk(clk));

lms_dsp_dspba_delay_10 d_u0_m0_wo0_wi0_r0_delayr15_q_11(
	.aclr(areset),
	.delay_signals_2_0(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][2]~q ),
	.delay_signals_9_0(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][9]~q ),
	.delay_signals_1_0(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][1]~q ),
	.delay_signals_8_0(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][8]~q ),
	.delay_signals_0_0(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][0]~q ),
	.delay_signals_7_0(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][3]~q ),
	.delay_signals_10_0(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][10]~q ),
	.delay_signals_11_0(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][11]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_43 u0_m0_wo0_wi0_r0_delayr15(
	.aclr(areset),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][2]~q ),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][9]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][1]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][8]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][0]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][3]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][0]~q }),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][10]~q ),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr15|delay_signals[0][11]~q ),
	.ena(xIn_v[0]),
	.clk(clk));

lms_dsp_dspba_delay_9 d_u0_m0_wo0_wi0_r0_delayr14_q_11(
	.aclr(areset),
	.delay_signals_4_0(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][2]~q ),
	.delay_signals_11_0(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][10]~q ),
	.delay_signals_9_0(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][5]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][2]~q ,gnd,gnd}),
	.clk(clk));

lms_dsp_dspba_delay_42 u0_m0_wo0_wi0_r0_delayr14(
	.aclr(areset),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][4]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][7]~q ),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][9]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][6]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][8]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][5]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][0]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][0]~q }),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][10]~q ),
	.ena(xIn_v[0]),
	.clk(clk));

lms_dsp_dspba_delay_8 d_u0_m0_wo0_wi0_r0_delayr13_q_11(
	.aclr(areset),
	.delay_signals_4_0(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][1]~q ),
	.delay_signals_11_0(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][10]~q ),
	.delay_signals_9_0(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][5]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][1]~q ,gnd}),
	.clk(clk));

lms_dsp_dspba_delay_41 u0_m0_wo0_wi0_r0_delayr13(
	.aclr(areset),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][4]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][6]~q ),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][9]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][5]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][7]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][0]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][0]~q }),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][10]~q ),
	.ena(xIn_v[0]),
	.clk(clk));

lms_dsp_dspba_delay_7 d_u0_m0_wo0_wi0_r0_delayr12_q_12(
	.aclr(areset),
	.delay_signals_6_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][1]~q ),
	.delay_signals_11_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][10]~q ),
	.delay_signals_9_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][7]~q ),
	.xin({\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][11]~q ,\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][10]~q ,\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][9]~q ,\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][8]~q ,
\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][7]~q ,\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][6]~q ,\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][5]~q ,\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][4]~q ,
\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][3]~q ,\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][2]~q ,\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][1]~q ,gnd}),
	.clk(clk));

lms_dsp_dspba_delay_6 d_u0_m0_wo0_wi0_r0_delayr12_q_11(
	.aclr(areset),
	.delay_signals_6_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][6]~q ),
	.delay_signals_8_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][8]~q ),
	.delay_signals_9_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][9]~q ),
	.delay_signals_7_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][7]~q ),
	.delay_signals_5_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][1]~q ),
	.delay_signals_0_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][0]~q ),
	.delay_signals_11_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][10]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_40 u0_m0_wo0_wi0_r0_delayr12(
	.aclr(areset),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][6]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][8]~q ),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][9]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][7]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][0]~q ),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr12|delay_signals[0][10]~q ),
	.ena(xIn_v[0]),
	.xin({\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_39 u0_m0_wo0_wi0_r0_delayr11(
	.aclr(areset),
	.xin({\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][0]~q }),
	.ena(xIn_v[0]),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][6]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][8]~q ),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][9]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][7]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][0]~q ),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr11|delay_signals[0][10]~q ),
	.clk(clk));

lms_dsp_dspba_delay_5 d_u0_m0_wo0_wi0_r0_delayr10_q_11(
	.aclr(areset),
	.delay_signals_7_0(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][1]~q ),
	.delay_signals_11_0(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][10]~q ),
	.delay_signals_9_0(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][8]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][1]~q ,gnd}),
	.clk(clk));

lms_dsp_dspba_delay_38 u0_m0_wo0_wi0_r0_delayr10(
	.aclr(areset),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][7]~q ),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][8]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][2]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][0]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][1]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][0]~q }),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][10]~q ),
	.ena(xIn_v[0]),
	.clk(clk));

lms_dsp_dspba_delay_20 d_u0_m0_wo0_wi0_r0_delayr9_q_11(
	.aclr(areset),
	.delay_signals_8_0(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][1]~q ),
	.delay_signals_0_0(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][0]~q ),
	.delay_signals_11_0(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][10]~q ),
	.delay_signals_9_0(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][9]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_61 u0_m0_wo0_wi0_r0_delayr9(
	.aclr(areset),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][0]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][0]~q }),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][10]~q ),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr9|delay_signals[0][9]~q ),
	.ena(xIn_v[0]),
	.clk(clk));

lms_dsp_dspba_delay_19 d_u0_m0_wo0_wi0_r0_delayr8_q_12(
	.aclr(areset),
	.delay_signals_7_0(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][7]~q ),
	.delay_signals_9_0(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][9]~q ),
	.delay_signals_6_0(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][6]~q ),
	.delay_signals_8_0(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][8]~q ),
	.delay_signals_5_0(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][1]~q ),
	.delay_signals_0_0(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][0]~q ),
	.delay_signals_10_0(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][10]~q ),
	.delay_signals_11_0(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][11]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_60 u0_m0_wo0_wi0_r0_delayr8(
	.aclr(areset),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][7]~q ),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][9]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][6]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][8]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][0]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][10]~q ),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr8|delay_signals[0][11]~q ),
	.ena(xIn_v[0]),
	.xin({\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_59 u0_m0_wo0_wi0_r0_delayr7(
	.aclr(areset),
	.xin({\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][0]~q }),
	.ena(xIn_v[0]),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][7]~q ),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][9]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][6]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][8]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][0]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][10]~q ),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr7|delay_signals[0][11]~q ),
	.clk(clk));

lms_dsp_dspba_delay_18 d_u0_m0_wo0_wi0_r0_delayr6_q_14(
	.aclr(areset),
	.delay_signals_9_0(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][1]~q ),
	.delay_signals_0_0(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][0]~q ),
	.delay_signals_11_0(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][10]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_58 u0_m0_wo0_wi0_r0_delayr6(
	.aclr(areset),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][9]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][0]~q }),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][0]~q ),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr6|delay_signals[0][10]~q ),
	.ena(xIn_v[0]),
	.clk(clk));

lms_dsp_dspba_delay_17 d_u0_m0_wo0_wi0_r0_delayr5_q_13(
	.aclr(areset),
	.delay_signals_9_0(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][2]~q ),
	.delay_signals_0_0(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][0]~q ),
	.delay_signals_1_0(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][1]~q ),
	.delay_signals_11_0(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][10]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_57 u0_m0_wo0_wi0_r0_delayr5(
	.aclr(areset),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][2]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][0]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][1]~q ),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr5|delay_signals[0][10]~q ),
	.ena(xIn_v[0]),
	.xin({\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_56 u0_m0_wo0_wi0_r0_delayr4(
	.aclr(areset),
	.ena(xIn_v[0]),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][2]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][0]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][1]~q ),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr4|delay_signals[0][10]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_55 u0_m0_wo0_wi0_r0_delayr3(
	.aclr(areset),
	.ena(xIn_v[0]),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][2]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][0]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][1]~q ),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr3|delay_signals[0][10]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_48 u0_m0_wo0_wi0_r0_delayr2(
	.aclr(areset),
	.ena(xIn_v[0]),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][2]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][0]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][1]~q ),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr2|delay_signals[0][10]~q ),
	.xin({\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][11]~q ,\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][10]~q ,\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][9]~q ,\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][8]~q ,\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][7]~q ,
\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][6]~q ,\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][5]~q ,\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][4]~q ,\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][3]~q ,\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][2]~q ,
\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][1]~q ,\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_37 u0_m0_wo0_wi0_r0_delayr1(
	.aclr(areset),
	.ena(xIn_v[0]),
	.delay_signals_9_0(\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][2]~q ),
	.delay_signals_0_0(\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][0]~q ),
	.delay_signals_1_0(\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][1]~q ),
	.delay_signals_11_0(\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u0_m0_wo0_wi0_r0_delayr1|delay_signals[0][10]~q ),
	.xin({xIn_0[11],xIn_0[10],xIn_0[9],xIn_0[8],xIn_0[7],xIn_0[6],xIn_0[5],xIn_0[4],xIn_0[3],xIn_0[2],xIn_0[1],xIn_0[0]}),
	.clk(clk));

lms_dsp_dspba_delay_79 u1_m0_wo0_wi0_r0_delayr25(
	.aclr(areset),
	.xin({\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][0]~q }),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][2]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][0]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][1]~q ),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][10]~q ),
	.ena(\d_u0_m0_wo0_compute_q_13|delay_signals[0][0]~q ),
	.clk(clk));

lms_dsp_dspba_delay_32 d_u1_m0_wo0_wi0_r0_delayr24_q_14(
	.aclr(areset),
	.delay_signals_9_0(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][1]~q ),
	.delay_signals_0_0(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][0]~q ),
	.delay_signals_11_0(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][10]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_78 u1_m0_wo0_wi0_r0_delayr24(
	.aclr(areset),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][0]~q ),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr24|delay_signals[0][10]~q ),
	.ena(\d_u0_m0_wo0_compute_q_13|delay_signals[0][0]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_77 u1_m0_wo0_wi0_r0_delayr23(
	.aclr(areset),
	.xin({\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][11]~q ,\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][10]~q ,\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][9]~q ,\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][8]~q ,
\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][7]~q ,\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][6]~q ,\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][5]~q ,\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][4]~q ,
\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][3]~q ,\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][2]~q ,\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][1]~q ,\u1_m0_wo0_mtree_add0_4_o[0]~q }),
	.ena(\d_u0_m0_wo0_compute_q_13|delay_signals[0][0]~q ),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][0]~q ),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr23|delay_signals[0][10]~q ),
	.clk(clk));

lms_dsp_dspba_delay_31 d_u1_m0_wo0_wi0_r0_delayr22_q_13(
	.aclr(areset),
	.u1_m0_wo0_mtree_mult1_8_sub_1_o_1(\u1_m0_wo0_mtree_mult1_8_sub_1_o[1]~q ),
	.delay_signals_9_0(\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][1]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][2]~q ,gnd,gnd}),
	.delay_signals_11_0(\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u1_m0_wo0_wi0_r0_delayr22_q_13|delay_signals[0][10]~q ),
	.clk(clk));

lms_dsp_dspba_delay_1 d_u0_m0_wo0_compute_q_13(
	.aclr(areset),
	.delay_signals_0_0(\d_u0_m0_wo0_compute_q_13|delay_signals[0][0]~q ),
	.xin({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\d_u0_m0_wo0_compute_q_11|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_76 u1_m0_wo0_wi0_r0_delayr22(
	.aclr(areset),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][7]~q ),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][9]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][6]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][8]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][0]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][0]~q }),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][10]~q ),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][11]~q ),
	.ena(\d_u0_m0_wo0_compute_q_11|delay_signals[0][0]~q ),
	.clk(clk));

lms_dsp_dspba_delay_75 u1_m0_wo0_wi0_r0_delayr21(
	.aclr(areset),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][0]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][0]~q }),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][10]~q ),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][9]~q ),
	.ena(\d_u0_m0_wo0_compute_q_11|delay_signals[0][0]~q ),
	.clk(clk));

lms_dsp_dspba_delay_30 d_u1_m0_wo0_wi0_r0_delayr20_q_12(
	.aclr(areset),
	.delay_signals_7_0(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][1]~q ),
	.delay_signals_11_0(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][10]~q ),
	.delay_signals_9_0(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][8]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][1]~q ,gnd}),
	.clk(clk));

lms_dsp_dspba_delay_74 u1_m0_wo0_wi0_r0_delayr20(
	.aclr(areset),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][7]~q ),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][8]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][2]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][0]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][1]~q ),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][10]~q ),
	.ena(\d_u0_m0_wo0_compute_q_11|delay_signals[0][0]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_72 u1_m0_wo0_wi0_r0_delayr19(
	.aclr(areset),
	.xin({\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][11]~q ,\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][10]~q ,\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][9]~q ,\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][8]~q ,
\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][7]~q ,\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][6]~q ,\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][5]~q ,\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][4]~q ,
\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][3]~q ,\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][2]~q ,\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][1]~q ,\u1_m0_wo0_mtree_mult1_12_add_1_o[0]~q }),
	.ena(\d_u0_m0_wo0_compute_q_11|delay_signals[0][0]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][7]~q ),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][8]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][2]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][0]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][1]~q ),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr19|delay_signals[0][10]~q ),
	.clk(clk));

lms_dsp_dspba_delay d_u0_m0_wo0_compute_q_11(
	.aclr(areset),
	.delay_signals_0_0(\d_u0_m0_wo0_compute_q_11|delay_signals[0][0]~q ),
	.xin({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,xIn_v[0]}),
	.clk(clk));

lms_dsp_dspba_delay_29 d_u1_m0_wo0_wi0_r0_delayr18_q_11(
	.aclr(areset),
	.delay_signals_6_0(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][1]~q ),
	.delay_signals_11_0(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][10]~q ),
	.delay_signals_9_0(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][7]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][1]~q ,gnd}),
	.clk(clk));

lms_dsp_dspba_delay_71 u1_m0_wo0_wi0_r0_delayr18(
	.aclr(areset),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][6]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][8]~q ),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][9]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][7]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][0]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][0]~q }),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][10]~q ),
	.ena(xIn_v[0]),
	.clk(clk));

lms_dsp_dspba_delay_28 d_u1_m0_wo0_wi0_r0_delayr17_q_11(
	.aclr(areset),
	.delay_signals_4_0(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][1]~q ),
	.delay_signals_11_0(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][10]~q ),
	.delay_signals_9_0(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][5]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][1]~q ,gnd}),
	.clk(clk));

lms_dsp_dspba_delay_70 u1_m0_wo0_wi0_r0_delayr17(
	.aclr(areset),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][4]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][6]~q ),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][9]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][5]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][7]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][0]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][0]~q }),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][10]~q ),
	.ena(xIn_v[0]),
	.clk(clk));

lms_dsp_dspba_delay_27 d_u1_m0_wo0_wi0_r0_delayr16_q_11(
	.aclr(areset),
	.delay_signals_4_0(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][2]~q ),
	.delay_signals_11_0(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][10]~q ),
	.delay_signals_9_0(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][5]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][2]~q ,gnd,gnd}),
	.clk(clk));

lms_dsp_dspba_delay_69 u1_m0_wo0_wi0_r0_delayr16(
	.aclr(areset),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][4]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][7]~q ),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][9]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][6]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][8]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][5]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][0]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][0]~q }),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][10]~q ),
	.ena(xIn_v[0]),
	.clk(clk));

lms_dsp_dspba_delay_26 d_u1_m0_wo0_wi0_r0_delayr15_q_11(
	.aclr(areset),
	.delay_signals_2_0(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][2]~q ),
	.delay_signals_9_0(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][9]~q ),
	.delay_signals_1_0(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][1]~q ),
	.delay_signals_8_0(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][8]~q ),
	.delay_signals_0_0(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][0]~q ),
	.delay_signals_7_0(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][3]~q ),
	.delay_signals_10_0(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][10]~q ),
	.delay_signals_11_0(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][11]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_68 u1_m0_wo0_wi0_r0_delayr15(
	.aclr(areset),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][2]~q ),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][9]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][1]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][8]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][0]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][3]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][0]~q }),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][10]~q ),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr15|delay_signals[0][11]~q ),
	.ena(xIn_v[0]),
	.clk(clk));

lms_dsp_dspba_delay_25 d_u1_m0_wo0_wi0_r0_delayr14_q_11(
	.aclr(areset),
	.delay_signals_4_0(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][2]~q ),
	.delay_signals_11_0(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][10]~q ),
	.delay_signals_9_0(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][5]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][2]~q ,gnd,gnd}),
	.clk(clk));

lms_dsp_dspba_delay_67 u1_m0_wo0_wi0_r0_delayr14(
	.aclr(areset),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][4]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][7]~q ),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][9]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][6]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][8]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][5]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][0]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][0]~q }),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][10]~q ),
	.ena(xIn_v[0]),
	.clk(clk));

lms_dsp_dspba_delay_24 d_u1_m0_wo0_wi0_r0_delayr13_q_11(
	.aclr(areset),
	.delay_signals_4_0(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][1]~q ),
	.delay_signals_11_0(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][10]~q ),
	.delay_signals_9_0(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][5]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][1]~q ,gnd}),
	.clk(clk));

lms_dsp_dspba_delay_66 u1_m0_wo0_wi0_r0_delayr13(
	.aclr(areset),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][4]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][6]~q ),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][9]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][5]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][7]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][0]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][0]~q }),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][10]~q ),
	.ena(xIn_v[0]),
	.clk(clk));

lms_dsp_dspba_delay_23 d_u1_m0_wo0_wi0_r0_delayr12_q_12(
	.aclr(areset),
	.delay_signals_6_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][1]~q ),
	.delay_signals_11_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][10]~q ),
	.delay_signals_9_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][7]~q ),
	.xin({\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][11]~q ,\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][10]~q ,\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][9]~q ,\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][8]~q ,
\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][7]~q ,\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][6]~q ,\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][5]~q ,\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][4]~q ,
\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][3]~q ,\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][2]~q ,\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][1]~q ,gnd}),
	.clk(clk));

lms_dsp_dspba_delay_22 d_u1_m0_wo0_wi0_r0_delayr12_q_11(
	.aclr(areset),
	.delay_signals_6_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][6]~q ),
	.delay_signals_8_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][8]~q ),
	.delay_signals_9_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][9]~q ),
	.delay_signals_7_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][7]~q ),
	.delay_signals_5_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][1]~q ),
	.delay_signals_0_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][0]~q ),
	.delay_signals_11_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][10]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_65 u1_m0_wo0_wi0_r0_delayr12(
	.aclr(areset),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][6]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][8]~q ),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][9]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][7]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][0]~q ),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr12|delay_signals[0][10]~q ),
	.ena(xIn_v[0]),
	.xin({\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_64 u1_m0_wo0_wi0_r0_delayr11(
	.aclr(areset),
	.xin({\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][0]~q }),
	.ena(xIn_v[0]),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][6]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][8]~q ),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][9]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][7]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][0]~q ),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr11|delay_signals[0][10]~q ),
	.clk(clk));

lms_dsp_dspba_delay_21 d_u1_m0_wo0_wi0_r0_delayr10_q_11(
	.aclr(areset),
	.delay_signals_7_0(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][1]~q ),
	.delay_signals_11_0(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][10]~q ),
	.delay_signals_9_0(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][8]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][1]~q ,gnd}),
	.clk(clk));

lms_dsp_dspba_delay_63 u1_m0_wo0_wi0_r0_delayr10(
	.aclr(areset),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][7]~q ),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][8]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][2]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][0]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][1]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][0]~q }),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][10]~q ),
	.ena(xIn_v[0]),
	.clk(clk));

lms_dsp_dspba_delay_36 d_u1_m0_wo0_wi0_r0_delayr9_q_11(
	.aclr(areset),
	.delay_signals_8_0(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][1]~q ),
	.delay_signals_0_0(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][0]~q ),
	.delay_signals_11_0(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][10]~q ),
	.delay_signals_9_0(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][9]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_86 u1_m0_wo0_wi0_r0_delayr9(
	.aclr(areset),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][0]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][0]~q }),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][10]~q ),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr9|delay_signals[0][9]~q ),
	.ena(xIn_v[0]),
	.clk(clk));

lms_dsp_dspba_delay_35 d_u1_m0_wo0_wi0_r0_delayr8_q_12(
	.aclr(areset),
	.delay_signals_7_0(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][7]~q ),
	.delay_signals_9_0(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][9]~q ),
	.delay_signals_6_0(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][6]~q ),
	.delay_signals_8_0(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][8]~q ),
	.delay_signals_5_0(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][1]~q ),
	.delay_signals_0_0(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][0]~q ),
	.delay_signals_10_0(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][10]~q ),
	.delay_signals_11_0(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][11]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_85 u1_m0_wo0_wi0_r0_delayr8(
	.aclr(areset),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][7]~q ),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][9]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][6]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][8]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][0]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][10]~q ),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr8|delay_signals[0][11]~q ),
	.ena(xIn_v[0]),
	.xin({\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_84 u1_m0_wo0_wi0_r0_delayr7(
	.aclr(areset),
	.xin({\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][0]~q }),
	.ena(xIn_v[0]),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][7]~q ),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][9]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][6]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][8]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][0]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][10]~q ),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr7|delay_signals[0][11]~q ),
	.clk(clk));

lms_dsp_dspba_delay_34 d_u1_m0_wo0_wi0_r0_delayr6_q_14(
	.aclr(areset),
	.delay_signals_9_0(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][2]~q ),
	.delay_signals_1_0(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][1]~q ),
	.delay_signals_0_0(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][0]~q ),
	.delay_signals_11_0(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][10]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_83 u1_m0_wo0_wi0_r0_delayr6(
	.aclr(areset),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][9]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][0]~q }),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][2]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][1]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][0]~q ),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr6|delay_signals[0][10]~q ),
	.ena(xIn_v[0]),
	.clk(clk));

lms_dsp_dspba_delay_33 d_u1_m0_wo0_wi0_r0_delayr5_q_13(
	.aclr(areset),
	.delay_signals_9_0(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][9]~q ),
	.delay_signals_8_0(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][8]~q ),
	.delay_signals_7_0(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][7]~q ),
	.delay_signals_6_0(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][6]~q ),
	.delay_signals_5_0(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][5]~q ),
	.delay_signals_4_0(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][4]~q ),
	.delay_signals_3_0(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][3]~q ),
	.delay_signals_2_0(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][2]~q ),
	.delay_signals_0_0(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][0]~q ),
	.delay_signals_1_0(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][1]~q ),
	.delay_signals_11_0(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][11]~q ),
	.delay_signals_10_0(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][10]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_82 u1_m0_wo0_wi0_r0_delayr5(
	.aclr(areset),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][2]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][0]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][1]~q ),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr5|delay_signals[0][10]~q ),
	.ena(xIn_v[0]),
	.xin({\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_81 u1_m0_wo0_wi0_r0_delayr4(
	.aclr(areset),
	.ena(xIn_v[0]),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][2]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][0]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][1]~q ),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr4|delay_signals[0][10]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_80 u1_m0_wo0_wi0_r0_delayr3(
	.aclr(areset),
	.ena(xIn_v[0]),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][2]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][0]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][1]~q ),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr3|delay_signals[0][10]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_73 u1_m0_wo0_wi0_r0_delayr2(
	.aclr(areset),
	.ena(xIn_v[0]),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][2]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][0]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][1]~q ),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr2|delay_signals[0][10]~q ),
	.xin({\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][11]~q ,\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][10]~q ,\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][9]~q ,\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][8]~q ,\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][7]~q ,
\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][6]~q ,\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][5]~q ,\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][4]~q ,\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][3]~q ,\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][2]~q ,
\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][1]~q ,\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][0]~q }),
	.clk(clk));

lms_dsp_dspba_delay_62 u1_m0_wo0_wi0_r0_delayr1(
	.aclr(areset),
	.ena(xIn_v[0]),
	.delay_signals_9_0(\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][9]~q ),
	.delay_signals_8_0(\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][8]~q ),
	.delay_signals_7_0(\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][7]~q ),
	.delay_signals_6_0(\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][6]~q ),
	.delay_signals_5_0(\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][5]~q ),
	.delay_signals_4_0(\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][4]~q ),
	.delay_signals_3_0(\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][3]~q ),
	.delay_signals_2_0(\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][2]~q ),
	.delay_signals_0_0(\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][0]~q ),
	.delay_signals_1_0(\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][1]~q ),
	.delay_signals_11_0(\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][11]~q ),
	.delay_signals_10_0(\u1_m0_wo0_wi0_r0_delayr1|delay_signals[0][10]~q ),
	.xin({xIn_1[11],xIn_1[10],xIn_1[9],xIn_1[8],xIn_1[7],xIn_1[6],xIn_1[5],xIn_1[4],xIn_1[3],xIn_1[2],xIn_1[1],xIn_1[0]}),
	.clk(clk));

dffeas \u1_m0_wo0_mtree_add4_0_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add4_0_o[9]~30_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u1_m0_wo0_mtree_add4_0_o_9),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add4_0_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add4_0_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add4_0_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add4_0_o[9]~30_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u0_m0_wo0_mtree_add4_0_o_9),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add4_0_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add4_0_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add4_0_o[20] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add4_0_o[20]~52_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u0_m0_wo0_mtree_add4_0_o_20),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add4_0_o[20] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add4_0_o[20] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add4_0_o[19] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add4_0_o[19]~50_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u0_m0_wo0_mtree_add4_0_o_19),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add4_0_o[19] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add4_0_o[19] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add4_0_o[18] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add4_0_o[18]~48_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u0_m0_wo0_mtree_add4_0_o_18),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add4_0_o[18] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add4_0_o[18] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add4_0_o[17] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add4_0_o[17]~46_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u0_m0_wo0_mtree_add4_0_o_17),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add4_0_o[17] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add4_0_o[17] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add4_0_o[16] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add4_0_o[16]~44_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u0_m0_wo0_mtree_add4_0_o_16),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add4_0_o[16] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add4_0_o[16] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add4_0_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add4_0_o[15]~42_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u0_m0_wo0_mtree_add4_0_o_15),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add4_0_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add4_0_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add4_0_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add4_0_o[14]~40_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u0_m0_wo0_mtree_add4_0_o_14),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add4_0_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add4_0_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add4_0_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add4_0_o[13]~38_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u0_m0_wo0_mtree_add4_0_o_13),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add4_0_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add4_0_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add4_0_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add4_0_o[12]~36_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u0_m0_wo0_mtree_add4_0_o_12),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add4_0_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add4_0_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add4_0_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add4_0_o[11]~34_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u0_m0_wo0_mtree_add4_0_o_11),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add4_0_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add4_0_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add4_0_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add4_0_o[10]~32_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u0_m0_wo0_mtree_add4_0_o_10),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add4_0_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add4_0_o[10] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add4_0_o[20] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add4_0_o[20]~52_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u1_m0_wo0_mtree_add4_0_o_20),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add4_0_o[20] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add4_0_o[20] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add4_0_o[19] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add4_0_o[19]~50_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u1_m0_wo0_mtree_add4_0_o_19),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add4_0_o[19] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add4_0_o[19] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add4_0_o[18] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add4_0_o[18]~48_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u1_m0_wo0_mtree_add4_0_o_18),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add4_0_o[18] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add4_0_o[18] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add4_0_o[17] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add4_0_o[17]~46_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u1_m0_wo0_mtree_add4_0_o_17),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add4_0_o[17] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add4_0_o[17] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add4_0_o[16] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add4_0_o[16]~44_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u1_m0_wo0_mtree_add4_0_o_16),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add4_0_o[16] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add4_0_o[16] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add4_0_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add4_0_o[15]~42_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u1_m0_wo0_mtree_add4_0_o_15),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add4_0_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add4_0_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add4_0_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add4_0_o[14]~40_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u1_m0_wo0_mtree_add4_0_o_14),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add4_0_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add4_0_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add4_0_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add4_0_o[13]~38_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u1_m0_wo0_mtree_add4_0_o_13),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add4_0_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add4_0_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add4_0_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add4_0_o[12]~36_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u1_m0_wo0_mtree_add4_0_o_12),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add4_0_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add4_0_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add4_0_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add4_0_o[11]~34_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u1_m0_wo0_mtree_add4_0_o_11),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add4_0_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add4_0_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add4_0_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add4_0_o[10]~32_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u1_m0_wo0_mtree_add4_0_o_10),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add4_0_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add4_0_o[10] .power_up = "low";

dffeas \u0_m0_wo0_oseq_gated_reg_q[0] (
	.clk(clk),
	.d(\d_u0_m0_wo0_compute_q_16|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(u0_m0_wo0_oseq_gated_reg_q_0),
	.prn(vcc));
defparam \u0_m0_wo0_oseq_gated_reg_q[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_oseq_gated_reg_q[0] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_5_sub_0_o[1]~12 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][0]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[1]~12_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[1]~13 ));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[1]~12 .lut_mask = 16'h6611;
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[1]~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_5_sub_0_o[2]~14 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_5_sub_0_o[1]~13 ),
	.combout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[2]~14_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[2]~15 ));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[2]~14 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[2]~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_5_sub_0_o[3]~16 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_5_sub_0_o[2]~15 ),
	.combout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[3]~16_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[3]~17 ));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[3]~16 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[3]~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_5_sub_0_o[4]~18 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_5_sub_0_o[3]~17 ),
	.combout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[4]~18_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[4]~19 ));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[4]~18 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[4]~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_5_sub_0_o[5]~20 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_5_sub_0_o[4]~19 ),
	.combout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[5]~20_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[5]~21 ));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[5]~20 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[5]~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_5_sub_0_o[6]~22 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_5_sub_0_o[5]~21 ),
	.combout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[6]~22_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[6]~23 ));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[6]~22 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[6]~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_5_sub_0_o[7]~24 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_5_sub_0_o[6]~23 ),
	.combout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[7]~24_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[7]~25 ));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[7]~24 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[7]~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_5_sub_0_o[8]~26 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_5_sub_0_o[7]~25 ),
	.combout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[8]~26_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[8]~27 ));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[8]~26 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[8]~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_5_sub_0_o[9]~28 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_5_sub_0_o[8]~27 ),
	.combout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[9]~28_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[9]~29 ));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[9]~28 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[9]~28 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_5_sub_0_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_5_sub_0_o[9]~28_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_5_sub_0_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_5_sub_0_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_5_sub_0_o[8]~26_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_5_sub_0_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_5_sub_0_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_5_sub_0_o[7]~24_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_5_sub_0_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_5_sub_0_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_5_sub_0_o[6]~22_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_5_sub_0_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_5_sub_0_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_5_sub_0_o[5]~20_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_5_sub_0_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_5_sub_0_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_5_sub_0_o[4]~18_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_5_sub_0_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_5_sub_0_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_5_sub_0_o[3]~16_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_5_sub_0_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_5_sub_0_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_5_sub_0_o[2]~14_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_5_sub_0_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_5_sub_0_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_5_sub_0_o[1]~12_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_5_sub_0_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_5_sub_0_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_5_sub_0_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_1_o[0]~14 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][0]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_5_sub_0_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_add1_1_o[0]~14_combout ),
	.cout(\u1_m0_wo0_mtree_add1_1_o[0]~15 ));
defparam \u1_m0_wo0_mtree_add1_1_o[0]~14 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_add1_1_o[0]~14 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_1_o[1]~16 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][1]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_5_sub_0_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_1_o[0]~15 ),
	.combout(\u1_m0_wo0_mtree_add1_1_o[1]~16_combout ),
	.cout(\u1_m0_wo0_mtree_add1_1_o[1]~17 ));
defparam \u1_m0_wo0_mtree_add1_1_o[1]~16 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_1_o[1]~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_1_o[2]~18 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][2]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_5_sub_0_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_1_o[1]~17 ),
	.combout(\u1_m0_wo0_mtree_add1_1_o[2]~18_combout ),
	.cout(\u1_m0_wo0_mtree_add1_1_o[2]~19 ));
defparam \u1_m0_wo0_mtree_add1_1_o[2]~18 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_1_o[2]~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_1_o[3]~20 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][3]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_5_sub_0_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_1_o[2]~19 ),
	.combout(\u1_m0_wo0_mtree_add1_1_o[3]~20_combout ),
	.cout(\u1_m0_wo0_mtree_add1_1_o[3]~21 ));
defparam \u1_m0_wo0_mtree_add1_1_o[3]~20 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_1_o[3]~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_1_o[4]~22 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][4]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_5_sub_0_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_1_o[3]~21 ),
	.combout(\u1_m0_wo0_mtree_add1_1_o[4]~22_combout ),
	.cout(\u1_m0_wo0_mtree_add1_1_o[4]~23 ));
defparam \u1_m0_wo0_mtree_add1_1_o[4]~22 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_1_o[4]~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_1_o[5]~24 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][5]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_5_sub_0_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_1_o[4]~23 ),
	.combout(\u1_m0_wo0_mtree_add1_1_o[5]~24_combout ),
	.cout(\u1_m0_wo0_mtree_add1_1_o[5]~25 ));
defparam \u1_m0_wo0_mtree_add1_1_o[5]~24 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_1_o[5]~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_1_o[6]~26 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][6]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_5_sub_0_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_1_o[5]~25 ),
	.combout(\u1_m0_wo0_mtree_add1_1_o[6]~26_combout ),
	.cout(\u1_m0_wo0_mtree_add1_1_o[6]~27 ));
defparam \u1_m0_wo0_mtree_add1_1_o[6]~26 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_1_o[6]~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_1_o[7]~28 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][7]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_5_sub_0_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_1_o[6]~27 ),
	.combout(\u1_m0_wo0_mtree_add1_1_o[7]~28_combout ),
	.cout(\u1_m0_wo0_mtree_add1_1_o[7]~29 ));
defparam \u1_m0_wo0_mtree_add1_1_o[7]~28 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_1_o[7]~28 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_1_o[8]~30 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][8]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_5_sub_0_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_1_o[7]~29 ),
	.combout(\u1_m0_wo0_mtree_add1_1_o[8]~30_combout ),
	.cout(\u1_m0_wo0_mtree_add1_1_o[8]~31 ));
defparam \u1_m0_wo0_mtree_add1_1_o[8]~30 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_1_o[8]~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_1_o[9]~32 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][9]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_5_sub_0_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_1_o[8]~31 ),
	.combout(\u1_m0_wo0_mtree_add1_1_o[9]~32_combout ),
	.cout(\u1_m0_wo0_mtree_add1_1_o[9]~33 ));
defparam \u1_m0_wo0_mtree_add1_1_o[9]~32 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_1_o[9]~32 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add1_1_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_1_o[9]~32_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_1_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_1_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_1_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_8_sub_1_o[2]~13 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][0]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[2]~13_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[2]~14 ));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[2]~13 .lut_mask = 16'h66DD;
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[2]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_8_sub_1_o[3]~15 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][1]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_8_sub_1_o[2]~14 ),
	.combout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[3]~15_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[3]~16 ));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[3]~15 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[3]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_8_sub_1_o[4]~17 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][2]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_8_sub_1_o[3]~16 ),
	.combout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[4]~17_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[4]~18 ));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[4]~17 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[4]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_8_sub_1_o[5]~19 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][3]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_8_sub_1_o[4]~18 ),
	.combout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[5]~19_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[5]~20 ));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[5]~19 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[5]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_8_sub_1_o[6]~21 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][4]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_8_sub_1_o[5]~20 ),
	.combout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[6]~21_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[6]~22 ));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[6]~21 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[6]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_8_sub_1_o[7]~23 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][5]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_8_sub_1_o[6]~22 ),
	.combout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[7]~23_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[7]~24 ));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[7]~23 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[7]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_8_sub_1_o[8]~25 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][6]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_8_sub_1_o[7]~24 ),
	.combout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[8]~25_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[8]~26 ));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[8]~25 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[8]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_8_sub_1_o[9]~27 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][7]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_8_sub_1_o[8]~26 ),
	.combout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[9]~27_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[9]~28 ));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[9]~27 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[9]~27 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_8_sub_1_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_8_sub_1_o[9]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_8_sub_1_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_9_add_1_o[1]~13 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][0]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_9_add_1_o[1]~13_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_9_add_1_o[1]~14 ));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[1]~13 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[1]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_9_add_1_o[2]~15 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][2]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_9_add_1_o[1]~14 ),
	.combout(\u1_m0_wo0_mtree_mult1_9_add_1_o[2]~15_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_9_add_1_o[2]~16 ));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[2]~15 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[2]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_9_add_1_o[3]~17 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][2]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_9_add_1_o[2]~16 ),
	.combout(\u1_m0_wo0_mtree_mult1_9_add_1_o[3]~17_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_9_add_1_o[3]~18 ));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[3]~17 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[3]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_9_add_1_o[4]~19 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][4]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_9_add_1_o[3]~18 ),
	.combout(\u1_m0_wo0_mtree_mult1_9_add_1_o[4]~19_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_9_add_1_o[4]~20 ));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[4]~19 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[4]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_9_add_1_o[5]~21 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][4]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_9_add_1_o[4]~20 ),
	.combout(\u1_m0_wo0_mtree_mult1_9_add_1_o[5]~21_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_9_add_1_o[5]~22 ));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[5]~21 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[5]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_9_add_1_o[6]~23 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][6]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_9_add_1_o[5]~22 ),
	.combout(\u1_m0_wo0_mtree_mult1_9_add_1_o[6]~23_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_9_add_1_o[6]~24 ));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[6]~23 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[6]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_9_add_1_o[7]~25 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][6]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_9_add_1_o[6]~24 ),
	.combout(\u1_m0_wo0_mtree_mult1_9_add_1_o[7]~25_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_9_add_1_o[7]~26 ));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[7]~25 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[7]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_9_add_1_o[8]~27 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][8]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_9_add_1_o[7]~26 ),
	.combout(\u1_m0_wo0_mtree_mult1_9_add_1_o[8]~27_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_9_add_1_o[8]~28 ));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[8]~27 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[8]~27 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_9_add_1_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_9_add_1_o[8]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_9_add_1_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_8_sub_1_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_8_sub_1_o[8]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_8_sub_1_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_9_add_1_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_9_add_1_o[7]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_9_add_1_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_8_sub_1_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_8_sub_1_o[7]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_8_sub_1_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_9_add_1_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_9_add_1_o[6]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_9_add_1_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_8_sub_1_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_8_sub_1_o[6]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_8_sub_1_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_9_add_1_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_9_add_1_o[5]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_9_add_1_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_8_sub_1_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_8_sub_1_o[5]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_8_sub_1_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_9_add_1_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_9_add_1_o[4]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_9_add_1_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_8_sub_1_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_8_sub_1_o[4]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_8_sub_1_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_9_add_1_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_9_add_1_o[3]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_9_add_1_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_8_sub_1_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_8_sub_1_o[3]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_8_sub_1_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_9_add_1_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_9_add_1_o[2]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_9_add_1_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_8_sub_1_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_8_sub_1_o[2]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_8_sub_1_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_9_add_1_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_9_add_1_o[1]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_9_add_1_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_8_sub_1_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_8_sub_1_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_9_add_1_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_9_add_1_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_4_o[1]~15 (
	.dataa(\u1_m0_wo0_mtree_mult1_8_sub_1_o[1]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_9_add_1_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_add0_4_o[1]~15_combout ),
	.cout(\u1_m0_wo0_mtree_add0_4_o[1]~16 ));
defparam \u1_m0_wo0_mtree_add0_4_o[1]~15 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_add0_4_o[1]~15 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_4_o[2]~17 (
	.dataa(\u1_m0_wo0_mtree_mult1_8_sub_1_o[2]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_9_add_1_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_4_o[1]~16 ),
	.combout(\u1_m0_wo0_mtree_add0_4_o[2]~17_combout ),
	.cout(\u1_m0_wo0_mtree_add0_4_o[2]~18 ));
defparam \u1_m0_wo0_mtree_add0_4_o[2]~17 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_4_o[2]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_4_o[3]~19 (
	.dataa(\u1_m0_wo0_mtree_mult1_8_sub_1_o[3]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_9_add_1_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_4_o[2]~18 ),
	.combout(\u1_m0_wo0_mtree_add0_4_o[3]~19_combout ),
	.cout(\u1_m0_wo0_mtree_add0_4_o[3]~20 ));
defparam \u1_m0_wo0_mtree_add0_4_o[3]~19 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_4_o[3]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_4_o[4]~21 (
	.dataa(\u1_m0_wo0_mtree_mult1_8_sub_1_o[4]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_9_add_1_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_4_o[3]~20 ),
	.combout(\u1_m0_wo0_mtree_add0_4_o[4]~21_combout ),
	.cout(\u1_m0_wo0_mtree_add0_4_o[4]~22 ));
defparam \u1_m0_wo0_mtree_add0_4_o[4]~21 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_4_o[4]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_4_o[5]~23 (
	.dataa(\u1_m0_wo0_mtree_mult1_8_sub_1_o[5]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_9_add_1_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_4_o[4]~22 ),
	.combout(\u1_m0_wo0_mtree_add0_4_o[5]~23_combout ),
	.cout(\u1_m0_wo0_mtree_add0_4_o[5]~24 ));
defparam \u1_m0_wo0_mtree_add0_4_o[5]~23 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_4_o[5]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_4_o[6]~25 (
	.dataa(\u1_m0_wo0_mtree_mult1_8_sub_1_o[6]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_9_add_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_4_o[5]~24 ),
	.combout(\u1_m0_wo0_mtree_add0_4_o[6]~25_combout ),
	.cout(\u1_m0_wo0_mtree_add0_4_o[6]~26 ));
defparam \u1_m0_wo0_mtree_add0_4_o[6]~25 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_4_o[6]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_4_o[7]~27 (
	.dataa(\u1_m0_wo0_mtree_mult1_8_sub_1_o[7]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_9_add_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_4_o[6]~26 ),
	.combout(\u1_m0_wo0_mtree_add0_4_o[7]~27_combout ),
	.cout(\u1_m0_wo0_mtree_add0_4_o[7]~28 ));
defparam \u1_m0_wo0_mtree_add0_4_o[7]~27 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_4_o[7]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_4_o[8]~29 (
	.dataa(\u1_m0_wo0_mtree_mult1_8_sub_1_o[8]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_9_add_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_4_o[7]~28 ),
	.combout(\u1_m0_wo0_mtree_add0_4_o[8]~29_combout ),
	.cout(\u1_m0_wo0_mtree_add0_4_o[8]~30 ));
defparam \u1_m0_wo0_mtree_add0_4_o[8]~29 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_4_o[8]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_4_o[9]~31 (
	.dataa(\u1_m0_wo0_mtree_mult1_8_sub_1_o[9]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_9_add_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_4_o[8]~30 ),
	.combout(\u1_m0_wo0_mtree_add0_4_o[9]~31_combout ),
	.cout(\u1_m0_wo0_mtree_add0_4_o[9]~32 ));
defparam \u1_m0_wo0_mtree_add0_4_o[9]~31 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_4_o[9]~31 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add0_4_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_4_o[9]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_4_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_4_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_4_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_0_o[1]~12 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][0]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[1]~12_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[1]~13 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[1]~12 .lut_mask = 16'h6611;
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[1]~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_0_o[2]~14 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_0_o[1]~13 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[2]~14_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[2]~15 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[2]~14 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[2]~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_0_o[3]~16 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_0_o[2]~15 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[3]~16_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[3]~17 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[3]~16 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[3]~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_0_o[4]~18 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_0_o[3]~17 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[4]~18_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[4]~19 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[4]~18 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[4]~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_0_o[5]~20 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_0_o[4]~19 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[5]~20_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[5]~21 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[5]~20 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[5]~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_0_o[6]~22 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_0_o[5]~21 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[6]~22_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[6]~23 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[6]~22 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[6]~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_0_o[7]~24 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_0_o[6]~23 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[7]~24_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[7]~25 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[7]~24 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[7]~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_0_o[8]~26 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_0_o[7]~25 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[8]~26_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[8]~27 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[8]~26 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[8]~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_0_o[9]~28 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_0_o[8]~27 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[9]~28_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[9]~29 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[9]~28 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[9]~28 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_0_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_0_o[9]~28_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_0_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_0_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_0_o[8]~26_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_0_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_0_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_0_o[7]~24_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_0_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_0_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_0_o[6]~22_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_0_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_0_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_0_o[5]~20_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_0_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_0_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_0_o[4]~18_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_0_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_0_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_0_o[3]~16_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_0_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_0_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_0_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_0_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_0_o[2]~14_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_0_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[2] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_2_o[2]~13 (
	.dataa(\u1_m0_wo0_mtree_mult1_10_sub_0_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_0_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[2]~13_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[2]~14 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[2]~13 .lut_mask = 16'h66DD;
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[2]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_2_o[3]~15 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][1]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_0_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_2_o[2]~14 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[3]~15_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[3]~16 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[3]~15 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[3]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_2_o[4]~17 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][2]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_0_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_2_o[3]~16 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[4]~17_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[4]~18 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[4]~17 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[4]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_2_o[5]~19 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][3]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_0_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_2_o[4]~18 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[5]~19_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[5]~20 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[5]~19 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[5]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_2_o[6]~21 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][4]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_0_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_2_o[5]~20 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[6]~21_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[6]~22 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[6]~21 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[6]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_2_o[7]~23 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][5]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_0_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_2_o[6]~22 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[7]~23_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[7]~24 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[7]~23 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[7]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_2_o[8]~25 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][6]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_0_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_2_o[7]~24 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[8]~25_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[8]~26 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[8]~25 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[8]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_2_o[9]~27 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][7]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_0_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_2_o[8]~26 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[9]~27_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[9]~28 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[9]~27 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[9]~27 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_2_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_2_o[9]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_2_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_4_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_4_o[8]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_4_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_4_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_4_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_2_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_2_o[8]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_2_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_4_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_4_o[7]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_4_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_4_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_4_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_2_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_2_o[7]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_2_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_4_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_4_o[6]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_4_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_4_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_4_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_2_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_2_o[6]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_2_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_4_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_4_o[5]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_4_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_4_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_4_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_2_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_2_o[5]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_2_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_4_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_4_o[4]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_4_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_4_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_4_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_2_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_2_o[4]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_2_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_4_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_4_o[3]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_4_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_4_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_4_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_2_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_2_o[3]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_2_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_4_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_4_o[2]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_4_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_4_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_4_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_2_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_2_o[2]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_2_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_4_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_4_o[1]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_4_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_4_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_4_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_0_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_0_o[1]~12_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_0_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_2_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_0_o[1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_2_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_8_sub_1_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_8_sub_1_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_4_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_8_sub_1_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_4_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_4_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_4_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_2_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_0_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_2_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_2_o[0]~17 (
	.dataa(\u1_m0_wo0_mtree_add0_4_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_2_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_add1_2_o[0]~17_combout ),
	.cout(\u1_m0_wo0_mtree_add1_2_o[0]~18 ));
defparam \u1_m0_wo0_mtree_add1_2_o[0]~17 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_add1_2_o[0]~17 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_2_o[1]~19 (
	.dataa(\u1_m0_wo0_mtree_add0_4_o[1]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_2_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_2_o[0]~18 ),
	.combout(\u1_m0_wo0_mtree_add1_2_o[1]~19_combout ),
	.cout(\u1_m0_wo0_mtree_add1_2_o[1]~20 ));
defparam \u1_m0_wo0_mtree_add1_2_o[1]~19 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_2_o[1]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_2_o[2]~21 (
	.dataa(\u1_m0_wo0_mtree_add0_4_o[2]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_2_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_2_o[1]~20 ),
	.combout(\u1_m0_wo0_mtree_add1_2_o[2]~21_combout ),
	.cout(\u1_m0_wo0_mtree_add1_2_o[2]~22 ));
defparam \u1_m0_wo0_mtree_add1_2_o[2]~21 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_2_o[2]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_2_o[3]~23 (
	.dataa(\u1_m0_wo0_mtree_add0_4_o[3]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_2_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_2_o[2]~22 ),
	.combout(\u1_m0_wo0_mtree_add1_2_o[3]~23_combout ),
	.cout(\u1_m0_wo0_mtree_add1_2_o[3]~24 ));
defparam \u1_m0_wo0_mtree_add1_2_o[3]~23 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_2_o[3]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_2_o[4]~25 (
	.dataa(\u1_m0_wo0_mtree_add0_4_o[4]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_2_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_2_o[3]~24 ),
	.combout(\u1_m0_wo0_mtree_add1_2_o[4]~25_combout ),
	.cout(\u1_m0_wo0_mtree_add1_2_o[4]~26 ));
defparam \u1_m0_wo0_mtree_add1_2_o[4]~25 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_2_o[4]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_2_o[5]~27 (
	.dataa(\u1_m0_wo0_mtree_add0_4_o[5]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_2_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_2_o[4]~26 ),
	.combout(\u1_m0_wo0_mtree_add1_2_o[5]~27_combout ),
	.cout(\u1_m0_wo0_mtree_add1_2_o[5]~28 ));
defparam \u1_m0_wo0_mtree_add1_2_o[5]~27 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_2_o[5]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_2_o[6]~29 (
	.dataa(\u1_m0_wo0_mtree_add0_4_o[6]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_2_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_2_o[5]~28 ),
	.combout(\u1_m0_wo0_mtree_add1_2_o[6]~29_combout ),
	.cout(\u1_m0_wo0_mtree_add1_2_o[6]~30 ));
defparam \u1_m0_wo0_mtree_add1_2_o[6]~29 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_2_o[6]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_2_o[7]~31 (
	.dataa(\u1_m0_wo0_mtree_add0_4_o[7]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_2_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_2_o[6]~30 ),
	.combout(\u1_m0_wo0_mtree_add1_2_o[7]~31_combout ),
	.cout(\u1_m0_wo0_mtree_add1_2_o[7]~32 ));
defparam \u1_m0_wo0_mtree_add1_2_o[7]~31 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_2_o[7]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_2_o[8]~33 (
	.dataa(\u1_m0_wo0_mtree_add0_4_o[8]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_2_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_2_o[7]~32 ),
	.combout(\u1_m0_wo0_mtree_add1_2_o[8]~33_combout ),
	.cout(\u1_m0_wo0_mtree_add1_2_o[8]~34 ));
defparam \u1_m0_wo0_mtree_add1_2_o[8]~33 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_2_o[8]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_2_o[9]~35 (
	.dataa(\u1_m0_wo0_mtree_add0_4_o[9]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_2_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_2_o[8]~34 ),
	.combout(\u1_m0_wo0_mtree_add1_2_o[9]~35_combout ),
	.cout(\u1_m0_wo0_mtree_add1_2_o[9]~36 ));
defparam \u1_m0_wo0_mtree_add1_2_o[9]~35 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_2_o[9]~35 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add1_2_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_2_o[9]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_2_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_2_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_2_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_1_o[1]~13 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][0]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_1_o[1]~13_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_1_o[1]~14 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[1]~13 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[1]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_1_o[2]~15 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][2]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_1_o[1]~14 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_1_o[2]~15_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_1_o[2]~16 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[2]~15 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[2]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_1_o[3]~17 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][2]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_1_o[2]~16 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_1_o[3]~17_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_1_o[3]~18 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[3]~17 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[3]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_1_o[4]~19 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][4]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_1_o[3]~18 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_1_o[4]~19_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_1_o[4]~20 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[4]~19 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[4]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_1_o[5]~21 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][4]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_1_o[4]~20 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_1_o[5]~21_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_1_o[5]~22 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[5]~21 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[5]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_1_o[6]~23 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][6]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_1_o[5]~22 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_1_o[6]~23_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_1_o[6]~24 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[6]~23 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[6]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_1_o[7]~25 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][6]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_1_o[6]~24 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_1_o[7]~25_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_1_o[7]~26 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[7]~25 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[7]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_1_o[8]~27 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][8]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_1_o[7]~26 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_1_o[8]~27_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_1_o[8]~28 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[8]~27 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[8]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_1_o[9]~29 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][8]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_1_o[8]~28 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_1_o[9]~29_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_1_o[9]~30 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[9]~29 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[9]~29 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_12_add_1_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_1_o[9]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_1_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_1_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_1_o[8]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_1_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_1_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_1_o[7]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_1_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_1_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_1_o[6]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_1_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_1_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_1_o[5]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_1_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_1_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_1_o[4]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_1_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_1_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_1_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_1_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_1_o[3]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_1_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[3] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_3_o[3]~13 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_1_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_12_add_1_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_3_o[3]~13_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_3_o[3]~14 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[3]~13 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[3]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_3_o[4]~15 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][1]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_12_add_1_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_3_o[3]~14 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_3_o[4]~15_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_3_o[4]~16 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[4]~15 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[4]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_3_o[5]~17 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][2]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_12_add_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_3_o[4]~16 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_3_o[5]~17_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_3_o[5]~18 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[5]~17 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[5]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_3_o[6]~19 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][3]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_12_add_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_3_o[5]~18 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_3_o[6]~19_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_3_o[6]~20 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[6]~19 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[6]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_3_o[7]~21 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][4]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_12_add_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_3_o[6]~20 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_3_o[7]~21_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_3_o[7]~22 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[7]~21 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[7]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_3_o[8]~23 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][5]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_12_add_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_3_o[7]~22 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_3_o[8]~23_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_3_o[8]~24 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[8]~23 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[8]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_3_o[9]~25 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][6]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_12_add_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_3_o[8]~24 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_3_o[9]~25_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_3_o[9]~26 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[9]~25 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[9]~25 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_12_add_3_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_3_o[9]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_3_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_1_o[1]~15 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][0]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[1]~15_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[1]~16 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[1]~15 .lut_mask = 16'h6611;
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[1]~15 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_1_o[2]~17 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_1_o[1]~16 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[2]~17_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[2]~18 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[2]~17 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[2]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_1_o[3]~19 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][0]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_1_o[2]~18 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[3]~19_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[3]~20 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[3]~19 .lut_mask = 16'h962B;
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[3]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_1_o[4]~21 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][1]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_1_o[3]~20 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[4]~21_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[4]~22 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[4]~21 .lut_mask = 16'h694D;
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[4]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_1_o[5]~23 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][2]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_1_o[4]~22 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[5]~23_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[5]~24 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[5]~23 .lut_mask = 16'h962B;
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[5]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_1_o[6]~25 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][3]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_1_o[5]~24 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[6]~25_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[6]~26 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[6]~25 .lut_mask = 16'h694D;
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[6]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_1_o[7]~27 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][4]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_1_o[6]~26 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[7]~27_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[7]~28 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[7]~27 .lut_mask = 16'h962B;
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[7]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_1_o[8]~29 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][5]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_1_o[7]~28 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[8]~29_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[8]~30 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[8]~29 .lut_mask = 16'h694D;
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[8]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_1_o[9]~31 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][6]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_1_o[8]~30 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[9]~31_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[9]~32 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[9]~31 .lut_mask = 16'h962B;
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[9]~31 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_1_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[9]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_1_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_1_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[8]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_1_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_1_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[7]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_1_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_1_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[6]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_1_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_1_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_1_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_1_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[5]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_1_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[5] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_3_o[5]~13 (
	.dataa(\u1_m0_wo0_mtree_mult1_13_sub_1_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[5]~13_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[5]~14 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[5]~13 .lut_mask = 16'h66DD;
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[5]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_3_o[6]~15 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][1]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_3_o[5]~14 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[6]~15_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[6]~16 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[6]~15 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[6]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_3_o[7]~17 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][2]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_3_o[6]~16 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[7]~17_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[7]~18 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[7]~17 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[7]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_3_o[8]~19 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][3]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_3_o[7]~18 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[8]~19_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[8]~20 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[8]~19 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[8]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_3_o[9]~21 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][4]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_3_o[8]~20 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[9]~21_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[9]~22 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[9]~21 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[9]~21 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_3_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_3_o[9]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_3_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_3_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_3_o[8]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_3_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_3_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_3_o[8]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_3_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_3_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_3_o[7]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_3_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_3_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_3_o[7]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_3_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_3_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_3_o[6]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_3_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_3_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_3_o[6]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_3_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_3_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_3_o[5]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_3_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_3_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_3_o[5]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_3_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_3_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_3_o[4]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_3_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_1_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[4]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_1_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_3_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[4]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_3_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_3_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_3_o[3]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_3_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_1_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[3]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_1_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_3_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[3]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_3_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_1_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_1_o[2]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_1_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_3_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_1_o[2]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_3_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_1_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[2]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_1_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_3_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[2]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_3_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_1_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_1_o[1]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_1_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_3_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_1_o[1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_3_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_1_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[1]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_1_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_3_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_3_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_3_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_1_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_3_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_3_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_3_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_6_o[0]~19 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_3_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_3_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_add0_6_o[0]~19_combout ),
	.cout(\u1_m0_wo0_mtree_add0_6_o[0]~20 ));
defparam \u1_m0_wo0_mtree_add0_6_o[0]~19 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_add0_6_o[0]~19 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_6_o[1]~21 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_3_o[1]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_3_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_6_o[0]~20 ),
	.combout(\u1_m0_wo0_mtree_add0_6_o[1]~21_combout ),
	.cout(\u1_m0_wo0_mtree_add0_6_o[1]~22 ));
defparam \u1_m0_wo0_mtree_add0_6_o[1]~21 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_6_o[1]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_6_o[2]~23 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_3_o[2]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_3_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_6_o[1]~22 ),
	.combout(\u1_m0_wo0_mtree_add0_6_o[2]~23_combout ),
	.cout(\u1_m0_wo0_mtree_add0_6_o[2]~24 ));
defparam \u1_m0_wo0_mtree_add0_6_o[2]~23 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_6_o[2]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_6_o[3]~25 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_3_o[3]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_3_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_6_o[2]~24 ),
	.combout(\u1_m0_wo0_mtree_add0_6_o[3]~25_combout ),
	.cout(\u1_m0_wo0_mtree_add0_6_o[3]~26 ));
defparam \u1_m0_wo0_mtree_add0_6_o[3]~25 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_6_o[3]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_6_o[4]~27 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_3_o[4]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_3_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_6_o[3]~26 ),
	.combout(\u1_m0_wo0_mtree_add0_6_o[4]~27_combout ),
	.cout(\u1_m0_wo0_mtree_add0_6_o[4]~28 ));
defparam \u1_m0_wo0_mtree_add0_6_o[4]~27 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_6_o[4]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_6_o[5]~29 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_3_o[5]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_3_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_6_o[4]~28 ),
	.combout(\u1_m0_wo0_mtree_add0_6_o[5]~29_combout ),
	.cout(\u1_m0_wo0_mtree_add0_6_o[5]~30 ));
defparam \u1_m0_wo0_mtree_add0_6_o[5]~29 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_6_o[5]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_6_o[6]~31 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_3_o[6]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_3_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_6_o[5]~30 ),
	.combout(\u1_m0_wo0_mtree_add0_6_o[6]~31_combout ),
	.cout(\u1_m0_wo0_mtree_add0_6_o[6]~32 ));
defparam \u1_m0_wo0_mtree_add0_6_o[6]~31 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_6_o[6]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_6_o[7]~33 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_3_o[7]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_3_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_6_o[6]~32 ),
	.combout(\u1_m0_wo0_mtree_add0_6_o[7]~33_combout ),
	.cout(\u1_m0_wo0_mtree_add0_6_o[7]~34 ));
defparam \u1_m0_wo0_mtree_add0_6_o[7]~33 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_6_o[7]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_6_o[8]~35 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_3_o[8]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_3_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_6_o[7]~34 ),
	.combout(\u1_m0_wo0_mtree_add0_6_o[8]~35_combout ),
	.cout(\u1_m0_wo0_mtree_add0_6_o[8]~36 ));
defparam \u1_m0_wo0_mtree_add0_6_o[8]~35 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_6_o[8]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_6_o[9]~37 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_3_o[9]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_3_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_6_o[8]~36 ),
	.combout(\u1_m0_wo0_mtree_add0_6_o[9]~37_combout ),
	.cout(\u1_m0_wo0_mtree_add0_6_o[9]~38 ));
defparam \u1_m0_wo0_mtree_add0_6_o[9]~37 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_6_o[9]~37 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add0_6_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_6_o[9]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_6_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_6_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_6_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_1_o[2]~13 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][0]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_1_o[2]~13_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_1_o[2]~14 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[2]~13 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[2]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_1_o[3]~15 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][1]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_1_o[2]~14 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_1_o[3]~15_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_1_o[3]~16 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[3]~15 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[3]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_1_o[4]~17 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][2]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_1_o[3]~16 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_1_o[4]~17_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_1_o[4]~18 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[4]~17 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[4]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_1_o[5]~19 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][3]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_1_o[4]~18 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_1_o[5]~19_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_1_o[5]~20 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[5]~19 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[5]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_1_o[6]~21 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][4]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_1_o[5]~20 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_1_o[6]~21_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_1_o[6]~22 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[6]~21 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[6]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_1_o[7]~23 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][5]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_1_o[6]~22 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_1_o[7]~23_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_1_o[7]~24 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[7]~23 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[7]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_1_o[8]~25 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][6]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_1_o[7]~24 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_1_o[8]~25_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_1_o[8]~26 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[8]~25 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[8]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_1_o[9]~27 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][7]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_1_o[8]~26 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_1_o[9]~27_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_1_o[9]~28 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[9]~27 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[9]~27 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_14_add_1_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_1_o[9]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_1_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_1_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_1_o[8]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_1_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_1_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_1_o[7]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_1_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_1_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_1_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_1_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_1_o[6]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_1_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_1_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_1_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_1_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_1_o[5]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_1_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[5] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_3_o[5]~13 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_1_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_14_add_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_3_o[5]~13_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_3_o[5]~14 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[5]~13 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[5]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_3_o[6]~15 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_1_o[1]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_14_add_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_3_o[5]~14 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_3_o[6]~15_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_3_o[6]~16 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[6]~15 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[6]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_3_o[7]~17 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][2]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_14_add_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_3_o[6]~16 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_3_o[7]~17_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_3_o[7]~18 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[7]~17 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[7]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_3_o[8]~19 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][3]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_14_add_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_3_o[7]~18 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_3_o[8]~19_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_3_o[8]~20 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[8]~19 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[8]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_3_o[9]~21 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][4]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_14_add_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_3_o[8]~20 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_3_o[9]~21_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_3_o[9]~22 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[9]~21 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[9]~21 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_14_add_3_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_3_o[9]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_3_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_15_sub_1_o[1]~19 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][0]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[1]~19_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[1]~20 ));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[1]~19 .lut_mask = 16'h6611;
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[1]~19 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_15_sub_1_o[2]~21 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_15_sub_1_o[1]~20 ),
	.combout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[2]~21_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[2]~22 ));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[2]~21 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[2]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_15_sub_1_o[3]~23 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_15_sub_1_o[2]~22 ),
	.combout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[3]~23_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[3]~24 ));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[3]~23 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[3]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_15_sub_1_o[4]~25 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_15_sub_1_o[3]~24 ),
	.combout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[4]~25_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[4]~26 ));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[4]~25 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[4]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_15_sub_1_o[5]~27 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_15_sub_1_o[4]~26 ),
	.combout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[5]~27_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[5]~28 ));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[5]~27 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[5]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_15_sub_1_o[6]~29 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_15_sub_1_o[5]~28 ),
	.combout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[6]~29_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[6]~30 ));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[6]~29 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[6]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_15_sub_1_o[7]~31 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][0]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_15_sub_1_o[6]~30 ),
	.combout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[7]~31_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[7]~32 ));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[7]~31 .lut_mask = 16'h962B;
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[7]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_15_sub_1_o[8]~33 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][1]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_15_sub_1_o[7]~32 ),
	.combout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[8]~33_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[8]~34 ));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[8]~33 .lut_mask = 16'h694D;
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[8]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_15_sub_1_o[9]~35 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][2]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_15_sub_1_o[8]~34 ),
	.combout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[9]~35_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[9]~36 ));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[9]~35 .lut_mask = 16'h962B;
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[9]~35 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_15_sub_1_o[9]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_3_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_3_o[8]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_3_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_15_sub_1_o[8]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_3_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_3_o[7]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_3_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_15_sub_1_o[7]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_3_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_3_o[6]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_3_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_15_sub_1_o[6]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_3_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_3_o[5]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_3_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_15_sub_1_o[5]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_1_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_1_o[4]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_1_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_3_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_1_o[4]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_3_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_15_sub_1_o[4]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_1_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_1_o[3]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_1_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_3_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_1_o[3]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_3_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_15_sub_1_o[3]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_1_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_1_o[2]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_1_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_3_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_1_o[2]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_3_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_15_sub_1_o[2]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_3_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_1_o[1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_3_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_15_sub_1_o[1]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_3_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_1_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_3_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[0] (
	.clk(clk),
	.d(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[0]~21 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_add0_7_o[0]~21_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[0]~22 ));
defparam \u1_m0_wo0_mtree_add0_7_o[0]~21 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_add0_7_o[0]~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[1]~23 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[1]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_7_o[0]~22 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[1]~23_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[1]~24 ));
defparam \u1_m0_wo0_mtree_add0_7_o[1]~23 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_7_o[1]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[2]~25 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[2]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_7_o[1]~24 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[2]~25_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[2]~26 ));
defparam \u1_m0_wo0_mtree_add0_7_o[2]~25 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_7_o[2]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[3]~27 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[3]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_7_o[2]~26 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[3]~27_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[3]~28 ));
defparam \u1_m0_wo0_mtree_add0_7_o[3]~27 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_7_o[3]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[4]~29 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[4]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_7_o[3]~28 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[4]~29_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[4]~30 ));
defparam \u1_m0_wo0_mtree_add0_7_o[4]~29 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_7_o[4]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[5]~31 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[5]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_7_o[4]~30 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[5]~31_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[5]~32 ));
defparam \u1_m0_wo0_mtree_add0_7_o[5]~31 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_7_o[5]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[6]~33 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[6]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_7_o[5]~32 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[6]~33_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[6]~34 ));
defparam \u1_m0_wo0_mtree_add0_7_o[6]~33 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_7_o[6]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[7]~35 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[7]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_7_o[6]~34 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[7]~35_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[7]~36 ));
defparam \u1_m0_wo0_mtree_add0_7_o[7]~35 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_7_o[7]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[8]~37 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[8]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_7_o[7]~36 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[8]~37_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[8]~38 ));
defparam \u1_m0_wo0_mtree_add0_7_o[8]~37 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_7_o[8]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[9]~39 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[9]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_7_o[8]~38 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[9]~39_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[9]~40 ));
defparam \u1_m0_wo0_mtree_add0_7_o[9]~39 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_7_o[9]~39 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add0_7_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[9]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_6_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_6_o[8]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_6_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_6_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_6_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_7_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[8]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_6_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_6_o[7]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_6_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_6_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_6_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_7_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[7]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_6_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_6_o[6]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_6_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_6_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_6_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_7_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[6]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_6_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_6_o[5]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_6_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_6_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_6_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_7_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[5]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_6_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_6_o[4]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_6_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_6_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_6_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_7_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[4]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_6_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_6_o[3]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_6_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_6_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_6_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_7_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[3]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_6_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_6_o[2]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_6_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_6_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_6_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_7_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[2]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_6_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_6_o[1]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_6_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_6_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_6_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_7_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[1]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_6_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_6_o[0]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_6_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_6_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_6_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_7_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[0]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[0]~21 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_add1_3_o[0]~21_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[0]~22 ));
defparam \u1_m0_wo0_mtree_add1_3_o[0]~21 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_add1_3_o[0]~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[1]~23 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[1]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_3_o[0]~22 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[1]~23_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[1]~24 ));
defparam \u1_m0_wo0_mtree_add1_3_o[1]~23 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_3_o[1]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[2]~25 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[2]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_3_o[1]~24 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[2]~25_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[2]~26 ));
defparam \u1_m0_wo0_mtree_add1_3_o[2]~25 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_3_o[2]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[3]~27 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[3]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_3_o[2]~26 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[3]~27_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[3]~28 ));
defparam \u1_m0_wo0_mtree_add1_3_o[3]~27 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_3_o[3]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[4]~29 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[4]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_3_o[3]~28 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[4]~29_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[4]~30 ));
defparam \u1_m0_wo0_mtree_add1_3_o[4]~29 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_3_o[4]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[5]~31 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[5]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_3_o[4]~30 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[5]~31_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[5]~32 ));
defparam \u1_m0_wo0_mtree_add1_3_o[5]~31 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_3_o[5]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[6]~33 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[6]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_3_o[5]~32 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[6]~33_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[6]~34 ));
defparam \u1_m0_wo0_mtree_add1_3_o[6]~33 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_3_o[6]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[7]~35 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[7]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_3_o[6]~34 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[7]~35_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[7]~36 ));
defparam \u1_m0_wo0_mtree_add1_3_o[7]~35 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_3_o[7]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[8]~37 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[8]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_3_o[7]~36 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[8]~37_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[8]~38 ));
defparam \u1_m0_wo0_mtree_add1_3_o[8]~37 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_3_o[8]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[9]~39 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[9]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_3_o[8]~38 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[9]~39_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[9]~40 ));
defparam \u1_m0_wo0_mtree_add1_3_o[9]~39 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_3_o[9]~39 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add1_3_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[9]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_2_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_2_o[8]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_2_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_2_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_2_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_3_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[8]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_2_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_2_o[7]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_2_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_2_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_2_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_3_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[7]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_2_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_2_o[6]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_2_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_2_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_2_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_3_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[6]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_2_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_2_o[5]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_2_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_2_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_2_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_3_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[5]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_2_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_2_o[4]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_2_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_2_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_2_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_3_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[4]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_2_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_2_o[3]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_2_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_2_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_2_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_3_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[3]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_2_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_2_o[2]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_2_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_2_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_2_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_3_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[2]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_2_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_2_o[1]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_2_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_2_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_2_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_3_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[1]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_2_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_2_o[0]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_2_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_2_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_2_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_3_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[0]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[0]~21 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_add2_1_o[0]~21_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[0]~22 ));
defparam \u1_m0_wo0_mtree_add2_1_o[0]~21 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_add2_1_o[0]~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[1]~23 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[1]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_1_o[0]~22 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[1]~23_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[1]~24 ));
defparam \u1_m0_wo0_mtree_add2_1_o[1]~23 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_1_o[1]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[2]~25 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[2]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_1_o[1]~24 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[2]~25_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[2]~26 ));
defparam \u1_m0_wo0_mtree_add2_1_o[2]~25 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add2_1_o[2]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[3]~27 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[3]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_1_o[2]~26 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[3]~27_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[3]~28 ));
defparam \u1_m0_wo0_mtree_add2_1_o[3]~27 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_1_o[3]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[4]~29 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[4]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_1_o[3]~28 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[4]~29_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[4]~30 ));
defparam \u1_m0_wo0_mtree_add2_1_o[4]~29 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add2_1_o[4]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[5]~31 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[5]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_1_o[4]~30 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[5]~31_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[5]~32 ));
defparam \u1_m0_wo0_mtree_add2_1_o[5]~31 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_1_o[5]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[6]~33 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[6]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_1_o[5]~32 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[6]~33_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[6]~34 ));
defparam \u1_m0_wo0_mtree_add2_1_o[6]~33 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add2_1_o[6]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[7]~35 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[7]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_1_o[6]~34 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[7]~35_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[7]~36 ));
defparam \u1_m0_wo0_mtree_add2_1_o[7]~35 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_1_o[7]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[8]~37 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[8]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_1_o[7]~36 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[8]~37_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[8]~38 ));
defparam \u1_m0_wo0_mtree_add2_1_o[8]~37 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add2_1_o[8]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[9]~39 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[9]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_1_o[8]~38 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[9]~39_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[9]~40 ));
defparam \u1_m0_wo0_mtree_add2_1_o[9]~39 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_1_o[9]~39 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add2_1_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[9]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_1_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_1_o[8]~30_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_1_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_1_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_1_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_1_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[8]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_1_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_1_o[7]~28_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_1_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_1_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_1_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_1_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[7]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_1_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_1_o[6]~26_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_1_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_1_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_1_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_1_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[6]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_1_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_1_o[5]~24_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_1_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_1_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_1_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_1_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[5]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_1_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_1_o[4]~22_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_1_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_1_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_1_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_1_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[4]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_1_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_1_o[3]~20_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_1_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_1_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_1_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_1_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[3]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_1_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_1_o[2]~18_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_1_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_1_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_1_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_1_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[2]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_1_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_1_o[1]~16_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_1_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_1_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_1_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_1_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[1]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_1_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_1_o[0]~14_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_1_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_1_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_1_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_1_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[0]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[0]~21 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_add3_0_o[0]~21_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[0]~22 ));
defparam \u1_m0_wo0_mtree_add3_0_o[0]~21 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_add3_0_o[0]~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[1]~23 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[1]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_0_o[0]~22 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[1]~23_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[1]~24 ));
defparam \u1_m0_wo0_mtree_add3_0_o[1]~23 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_0_o[1]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[2]~25 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[2]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_0_o[1]~24 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[2]~25_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[2]~26 ));
defparam \u1_m0_wo0_mtree_add3_0_o[2]~25 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add3_0_o[2]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[3]~27 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[3]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_0_o[2]~26 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[3]~27_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[3]~28 ));
defparam \u1_m0_wo0_mtree_add3_0_o[3]~27 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_0_o[3]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[4]~29 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[4]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_0_o[3]~28 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[4]~29_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[4]~30 ));
defparam \u1_m0_wo0_mtree_add3_0_o[4]~29 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add3_0_o[4]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[5]~31 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[5]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_0_o[4]~30 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[5]~31_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[5]~32 ));
defparam \u1_m0_wo0_mtree_add3_0_o[5]~31 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_0_o[5]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[6]~33 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[6]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_0_o[5]~32 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[6]~33_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[6]~34 ));
defparam \u1_m0_wo0_mtree_add3_0_o[6]~33 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add3_0_o[6]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[7]~35 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[7]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_0_o[6]~34 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[7]~35_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[7]~36 ));
defparam \u1_m0_wo0_mtree_add3_0_o[7]~35 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_0_o[7]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[8]~37 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[8]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_0_o[7]~36 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[8]~37_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[8]~38 ));
defparam \u1_m0_wo0_mtree_add3_0_o[8]~37 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add3_0_o[8]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[9]~39 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[9]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_0_o[8]~38 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[9]~39_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[9]~40 ));
defparam \u1_m0_wo0_mtree_add3_0_o[9]~39 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_0_o[9]~39 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add3_0_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[9]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_1_o[2]~13 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][0]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_1_o[2]~13_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_1_o[2]~14 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[2]~13 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[2]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_1_o[3]~15 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][1]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_1_o[2]~14 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_1_o[3]~15_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_1_o[3]~16 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[3]~15 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[3]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_1_o[4]~17 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][2]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_1_o[3]~16 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_1_o[4]~17_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_1_o[4]~18 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[4]~17 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[4]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_1_o[5]~19 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][3]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_1_o[4]~18 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_1_o[5]~19_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_1_o[5]~20 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[5]~19 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[5]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_1_o[6]~21 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][4]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_1_o[5]~20 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_1_o[6]~21_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_1_o[6]~22 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[6]~21 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[6]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_1_o[7]~23 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][5]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_1_o[6]~22 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_1_o[7]~23_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_1_o[7]~24 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[7]~23 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[7]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_1_o[8]~25 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][6]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_1_o[7]~24 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_1_o[8]~25_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_1_o[8]~26 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[8]~25 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[8]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_1_o[9]~27 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][7]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_1_o[8]~26 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_1_o[9]~27_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_1_o[9]~28 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[9]~27 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[9]~27 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_16_add_1_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_1_o[9]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_1_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_1_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_1_o[8]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_1_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_1_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_1_o[7]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_1_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_1_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_1_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_1_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_1_o[6]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_1_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_1_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_1_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_1_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_1_o[5]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_1_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[5] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_3_o[5]~13 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_1_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_16_add_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_3_o[5]~13_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_3_o[5]~14 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[5]~13 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[5]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_3_o[6]~15 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_1_o[1]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_16_add_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_3_o[5]~14 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_3_o[6]~15_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_3_o[6]~16 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[6]~15 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[6]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_3_o[7]~17 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][2]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_16_add_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_3_o[6]~16 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_3_o[7]~17_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_3_o[7]~18 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[7]~17 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[7]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_3_o[8]~19 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][3]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_16_add_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_3_o[7]~18 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_3_o[8]~19_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_3_o[8]~20 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[8]~19 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[8]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_3_o[9]~21 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][4]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_16_add_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_3_o[8]~20 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_3_o[9]~21_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_3_o[9]~22 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[9]~21 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[9]~21 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_16_add_3_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_3_o[9]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_3_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_1_o[1]~15 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][0]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[1]~15_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[1]~16 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[1]~15 .lut_mask = 16'h6611;
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[1]~15 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_1_o[2]~17 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_1_o[1]~16 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[2]~17_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[2]~18 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[2]~17 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[2]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_1_o[3]~19 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][0]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_1_o[2]~18 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[3]~19_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[3]~20 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[3]~19 .lut_mask = 16'h962B;
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[3]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_1_o[4]~21 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][1]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_1_o[3]~20 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[4]~21_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[4]~22 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[4]~21 .lut_mask = 16'h694D;
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[4]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_1_o[5]~23 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][2]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_1_o[4]~22 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[5]~23_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[5]~24 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[5]~23 .lut_mask = 16'h962B;
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[5]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_1_o[6]~25 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][3]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_1_o[5]~24 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[6]~25_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[6]~26 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[6]~25 .lut_mask = 16'h694D;
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[6]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_1_o[7]~27 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][4]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_1_o[6]~26 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[7]~27_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[7]~28 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[7]~27 .lut_mask = 16'h962B;
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[7]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_1_o[8]~29 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][5]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_1_o[7]~28 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[8]~29_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[8]~30 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[8]~29 .lut_mask = 16'h694D;
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[8]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_1_o[9]~31 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][6]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_1_o[8]~30 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[9]~31_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[9]~32 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[9]~31 .lut_mask = 16'h962B;
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[9]~31 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_1_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[9]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_1_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_1_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[8]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_1_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_1_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[7]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_1_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_1_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[6]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_1_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_1_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_1_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_1_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[5]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_1_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[5] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_3_o[5]~13 (
	.dataa(\u1_m0_wo0_mtree_mult1_17_sub_1_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[5]~13_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[5]~14 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[5]~13 .lut_mask = 16'h66DD;
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[5]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_3_o[6]~15 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][1]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_3_o[5]~14 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[6]~15_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[6]~16 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[6]~15 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[6]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_3_o[7]~17 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][2]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_3_o[6]~16 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[7]~17_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[7]~18 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[7]~17 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[7]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_3_o[8]~19 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][3]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_3_o[7]~18 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[8]~19_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[8]~20 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[8]~19 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[8]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_3_o[9]~21 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][4]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_3_o[8]~20 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[9]~21_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[9]~22 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[9]~21 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[9]~21 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_3_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_3_o[9]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_3_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_3_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_3_o[8]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_3_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_3_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_3_o[8]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_3_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_3_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_3_o[7]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_3_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_3_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_3_o[7]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_3_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_3_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_3_o[6]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_3_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_3_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_3_o[6]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_3_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_3_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_3_o[5]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_3_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_3_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_3_o[5]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_3_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_1_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_1_o[4]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_1_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_3_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_1_o[4]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_3_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_1_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[4]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_1_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_3_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[4]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_3_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_1_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_1_o[3]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_1_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_3_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_1_o[3]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_3_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_1_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[3]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_1_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_3_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[3]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_3_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_1_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_1_o[2]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_1_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_3_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_1_o[2]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_3_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_1_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[2]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_1_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_3_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[2]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_3_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_3_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_1_o[1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_3_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_1_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[1]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_1_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_3_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_3_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_3_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_1_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_3_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_3_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_3_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_8_o[0]~19 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_3_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_3_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_add0_8_o[0]~19_combout ),
	.cout(\u1_m0_wo0_mtree_add0_8_o[0]~20 ));
defparam \u1_m0_wo0_mtree_add0_8_o[0]~19 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_add0_8_o[0]~19 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_8_o[1]~21 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_3_o[1]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_3_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_8_o[0]~20 ),
	.combout(\u1_m0_wo0_mtree_add0_8_o[1]~21_combout ),
	.cout(\u1_m0_wo0_mtree_add0_8_o[1]~22 ));
defparam \u1_m0_wo0_mtree_add0_8_o[1]~21 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_8_o[1]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_8_o[2]~23 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_3_o[2]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_3_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_8_o[1]~22 ),
	.combout(\u1_m0_wo0_mtree_add0_8_o[2]~23_combout ),
	.cout(\u1_m0_wo0_mtree_add0_8_o[2]~24 ));
defparam \u1_m0_wo0_mtree_add0_8_o[2]~23 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_8_o[2]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_8_o[3]~25 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_3_o[3]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_3_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_8_o[2]~24 ),
	.combout(\u1_m0_wo0_mtree_add0_8_o[3]~25_combout ),
	.cout(\u1_m0_wo0_mtree_add0_8_o[3]~26 ));
defparam \u1_m0_wo0_mtree_add0_8_o[3]~25 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_8_o[3]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_8_o[4]~27 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_3_o[4]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_3_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_8_o[3]~26 ),
	.combout(\u1_m0_wo0_mtree_add0_8_o[4]~27_combout ),
	.cout(\u1_m0_wo0_mtree_add0_8_o[4]~28 ));
defparam \u1_m0_wo0_mtree_add0_8_o[4]~27 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_8_o[4]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_8_o[5]~29 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_3_o[5]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_3_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_8_o[4]~28 ),
	.combout(\u1_m0_wo0_mtree_add0_8_o[5]~29_combout ),
	.cout(\u1_m0_wo0_mtree_add0_8_o[5]~30 ));
defparam \u1_m0_wo0_mtree_add0_8_o[5]~29 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_8_o[5]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_8_o[6]~31 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_3_o[6]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_3_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_8_o[5]~30 ),
	.combout(\u1_m0_wo0_mtree_add0_8_o[6]~31_combout ),
	.cout(\u1_m0_wo0_mtree_add0_8_o[6]~32 ));
defparam \u1_m0_wo0_mtree_add0_8_o[6]~31 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_8_o[6]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_8_o[7]~33 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_3_o[7]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_3_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_8_o[6]~32 ),
	.combout(\u1_m0_wo0_mtree_add0_8_o[7]~33_combout ),
	.cout(\u1_m0_wo0_mtree_add0_8_o[7]~34 ));
defparam \u1_m0_wo0_mtree_add0_8_o[7]~33 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_8_o[7]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_8_o[8]~35 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_3_o[8]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_3_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_8_o[7]~34 ),
	.combout(\u1_m0_wo0_mtree_add0_8_o[8]~35_combout ),
	.cout(\u1_m0_wo0_mtree_add0_8_o[8]~36 ));
defparam \u1_m0_wo0_mtree_add0_8_o[8]~35 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_8_o[8]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_8_o[9]~37 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_3_o[9]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_3_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_8_o[8]~36 ),
	.combout(\u1_m0_wo0_mtree_add0_8_o[9]~37_combout ),
	.cout(\u1_m0_wo0_mtree_add0_8_o[9]~38 ));
defparam \u1_m0_wo0_mtree_add0_8_o[9]~37 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_8_o[9]~37 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add0_8_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_8_o[9]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_8_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_8_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_8_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_1_o[1]~13 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][0]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_1_o[1]~13_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_1_o[1]~14 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[1]~13 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[1]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_1_o[2]~15 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][2]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_1_o[1]~14 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_1_o[2]~15_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_1_o[2]~16 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[2]~15 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[2]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_1_o[3]~17 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][2]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_1_o[2]~16 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_1_o[3]~17_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_1_o[3]~18 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[3]~17 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[3]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_1_o[4]~19 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][4]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_1_o[3]~18 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_1_o[4]~19_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_1_o[4]~20 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[4]~19 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[4]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_1_o[5]~21 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][4]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_1_o[4]~20 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_1_o[5]~21_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_1_o[5]~22 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[5]~21 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[5]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_1_o[6]~23 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][6]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_1_o[5]~22 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_1_o[6]~23_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_1_o[6]~24 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[6]~23 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[6]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_1_o[7]~25 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][6]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_1_o[6]~24 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_1_o[7]~25_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_1_o[7]~26 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[7]~25 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[7]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_1_o[8]~27 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][8]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_1_o[7]~26 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_1_o[8]~27_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_1_o[8]~28 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[8]~27 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[8]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_1_o[9]~29 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][8]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_1_o[8]~28 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_1_o[9]~29_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_1_o[9]~30 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[9]~29 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[9]~29 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_18_add_1_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_1_o[9]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_1_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_1_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_1_o[8]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_1_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_1_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_1_o[7]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_1_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_1_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_1_o[6]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_1_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_1_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_1_o[5]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_1_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_1_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_1_o[4]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_1_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_1_o[0] (
	.clk(clk),
	.d(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_1_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_1_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_1_o[3]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_1_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[3] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_3_o[3]~13 (
	.dataa(\u1_m0_wo0_mtree_mult1_18_add_1_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_1_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_3_o[3]~13_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_3_o[3]~14 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[3]~13 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[3]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_3_o[4]~15 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][1]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_1_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_3_o[3]~14 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_3_o[4]~15_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_3_o[4]~16 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[4]~15 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[4]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_3_o[5]~17 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][2]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_3_o[4]~16 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_3_o[5]~17_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_3_o[5]~18 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[5]~17 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[5]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_3_o[6]~19 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][3]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_3_o[5]~18 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_3_o[6]~19_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_3_o[6]~20 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[6]~19 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[6]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_3_o[7]~21 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][4]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_3_o[6]~20 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_3_o[7]~21_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_3_o[7]~22 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[7]~21 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[7]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_3_o[8]~23 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][5]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_3_o[7]~22 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_3_o[8]~23_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_3_o[8]~24 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[8]~23 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[8]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_3_o[9]~25 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][6]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_3_o[8]~24 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_3_o[9]~25_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_3_o[9]~26 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[9]~25 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[9]~25 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_18_add_3_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_3_o[9]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_3_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_8_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_8_o[8]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_8_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_8_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_8_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_3_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_3_o[8]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_3_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_8_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_8_o[7]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_8_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_8_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_8_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_3_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_3_o[7]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_3_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_8_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_8_o[6]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_8_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_8_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_8_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_3_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_3_o[6]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_3_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_8_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_8_o[5]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_8_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_8_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_8_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_3_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_3_o[5]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_3_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_8_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_8_o[4]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_8_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_8_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_8_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_3_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_3_o[4]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_3_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_8_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_8_o[3]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_8_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_8_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_8_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_3_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_3_o[3]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_3_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_8_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_8_o[2]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_8_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_8_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_8_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_1_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_1_o[2]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_1_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_3_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_1_o[2]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_3_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_8_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_8_o[1]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_8_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_8_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_8_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_1_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_1_o[1]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_1_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_3_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_1_o[1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_3_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_8_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_8_o[0]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_8_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_8_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_8_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_3_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_1_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_3_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[0]~20 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_add1_4_o[0]~20_combout ),
	.cout(\u1_m0_wo0_mtree_add1_4_o[0]~21 ));
defparam \u1_m0_wo0_mtree_add1_4_o[0]~20 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_add1_4_o[0]~20 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[1]~22 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[1]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_4_o[0]~21 ),
	.combout(\u1_m0_wo0_mtree_add1_4_o[1]~22_combout ),
	.cout(\u1_m0_wo0_mtree_add1_4_o[1]~23 ));
defparam \u1_m0_wo0_mtree_add1_4_o[1]~22 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_4_o[1]~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[2]~24 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[2]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_4_o[1]~23 ),
	.combout(\u1_m0_wo0_mtree_add1_4_o[2]~24_combout ),
	.cout(\u1_m0_wo0_mtree_add1_4_o[2]~25 ));
defparam \u1_m0_wo0_mtree_add1_4_o[2]~24 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_4_o[2]~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[3]~26 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[3]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_4_o[2]~25 ),
	.combout(\u1_m0_wo0_mtree_add1_4_o[3]~26_combout ),
	.cout(\u1_m0_wo0_mtree_add1_4_o[3]~27 ));
defparam \u1_m0_wo0_mtree_add1_4_o[3]~26 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_4_o[3]~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[4]~28 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[4]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_4_o[3]~27 ),
	.combout(\u1_m0_wo0_mtree_add1_4_o[4]~28_combout ),
	.cout(\u1_m0_wo0_mtree_add1_4_o[4]~29 ));
defparam \u1_m0_wo0_mtree_add1_4_o[4]~28 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_4_o[4]~28 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[5]~30 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[5]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_4_o[4]~29 ),
	.combout(\u1_m0_wo0_mtree_add1_4_o[5]~30_combout ),
	.cout(\u1_m0_wo0_mtree_add1_4_o[5]~31 ));
defparam \u1_m0_wo0_mtree_add1_4_o[5]~30 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_4_o[5]~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[6]~32 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[6]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_4_o[5]~31 ),
	.combout(\u1_m0_wo0_mtree_add1_4_o[6]~32_combout ),
	.cout(\u1_m0_wo0_mtree_add1_4_o[6]~33 ));
defparam \u1_m0_wo0_mtree_add1_4_o[6]~32 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_4_o[6]~32 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[7]~34 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[7]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_4_o[6]~33 ),
	.combout(\u1_m0_wo0_mtree_add1_4_o[7]~34_combout ),
	.cout(\u1_m0_wo0_mtree_add1_4_o[7]~35 ));
defparam \u1_m0_wo0_mtree_add1_4_o[7]~34 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_4_o[7]~34 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[8]~36 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[8]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_4_o[7]~35 ),
	.combout(\u1_m0_wo0_mtree_add1_4_o[8]~36_combout ),
	.cout(\u1_m0_wo0_mtree_add1_4_o[8]~37 ));
defparam \u1_m0_wo0_mtree_add1_4_o[8]~36 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_4_o[8]~36 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[9]~38 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[9]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_4_o[8]~37 ),
	.combout(\u1_m0_wo0_mtree_add1_4_o[9]~38_combout ),
	.cout(\u1_m0_wo0_mtree_add1_4_o[9]~39 ));
defparam \u1_m0_wo0_mtree_add1_4_o[9]~38 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_4_o[9]~38 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add1_4_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[9]~38_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_0_o[1]~12 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][0]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[1]~12_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[1]~13 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[1]~12 .lut_mask = 16'h6611;
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[1]~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_0_o[2]~14 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_0_o[1]~13 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[2]~14_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[2]~15 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[2]~14 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[2]~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_0_o[3]~16 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_0_o[2]~15 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[3]~16_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[3]~17 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[3]~16 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[3]~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_0_o[4]~18 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_0_o[3]~17 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[4]~18_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[4]~19 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[4]~18 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[4]~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_0_o[5]~20 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_0_o[4]~19 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[5]~20_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[5]~21 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[5]~20 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[5]~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_0_o[6]~22 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_0_o[5]~21 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[6]~22_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[6]~23 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[6]~22 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[6]~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_0_o[7]~24 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_0_o[6]~23 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[7]~24_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[7]~25 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[7]~24 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[7]~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_0_o[8]~26 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_0_o[7]~25 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[8]~26_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[8]~27 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[8]~26 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[8]~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_0_o[9]~28 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_0_o[8]~27 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[9]~28_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[9]~29 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[9]~28 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[9]~28 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_0_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_0_o[9]~28_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_0_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_0_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_0_o[8]~26_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_0_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_0_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_0_o[7]~24_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_0_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_0_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_0_o[6]~22_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_0_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_0_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_0_o[5]~20_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_0_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_0_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_0_o[4]~18_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_0_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_0_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_0_o[3]~16_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_0_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_0_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_0_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_0_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_0_o[2]~14_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_0_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[2] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_2_o[2]~13 (
	.dataa(\u1_m0_wo0_mtree_mult1_20_sub_0_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_20_sub_0_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[2]~13_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[2]~14 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[2]~13 .lut_mask = 16'h66DD;
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[2]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_2_o[3]~15 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][1]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_20_sub_0_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_2_o[2]~14 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[3]~15_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[3]~16 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[3]~15 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[3]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_2_o[4]~17 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][2]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_20_sub_0_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_2_o[3]~16 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[4]~17_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[4]~18 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[4]~17 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[4]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_2_o[5]~19 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][3]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_20_sub_0_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_2_o[4]~18 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[5]~19_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[5]~20 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[5]~19 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[5]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_2_o[6]~21 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][4]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_20_sub_0_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_2_o[5]~20 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[6]~21_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[6]~22 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[6]~21 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[6]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_2_o[7]~23 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][5]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_20_sub_0_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_2_o[6]~22 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[7]~23_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[7]~24 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[7]~23 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[7]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_2_o[8]~25 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][6]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_20_sub_0_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_2_o[7]~24 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[8]~25_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[8]~26 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[8]~25 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[8]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_2_o[9]~27 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][7]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_20_sub_0_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_2_o[8]~26 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[9]~27_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[9]~28 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[9]~27 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[9]~27 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_2_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_2_o[9]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_2_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_21_add_1_o[1]~13 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][0]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_21_add_1_o[1]~13_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_21_add_1_o[1]~14 ));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[1]~13 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[1]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_21_add_1_o[2]~15 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][2]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_21_add_1_o[1]~14 ),
	.combout(\u1_m0_wo0_mtree_mult1_21_add_1_o[2]~15_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_21_add_1_o[2]~16 ));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[2]~15 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[2]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_21_add_1_o[3]~17 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][2]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_21_add_1_o[2]~16 ),
	.combout(\u1_m0_wo0_mtree_mult1_21_add_1_o[3]~17_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_21_add_1_o[3]~18 ));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[3]~17 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[3]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_21_add_1_o[4]~19 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][4]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_21_add_1_o[3]~18 ),
	.combout(\u1_m0_wo0_mtree_mult1_21_add_1_o[4]~19_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_21_add_1_o[4]~20 ));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[4]~19 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[4]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_21_add_1_o[5]~21 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][4]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_21_add_1_o[4]~20 ),
	.combout(\u1_m0_wo0_mtree_mult1_21_add_1_o[5]~21_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_21_add_1_o[5]~22 ));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[5]~21 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[5]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_21_add_1_o[6]~23 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][6]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_21_add_1_o[5]~22 ),
	.combout(\u1_m0_wo0_mtree_mult1_21_add_1_o[6]~23_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_21_add_1_o[6]~24 ));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[6]~23 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[6]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_21_add_1_o[7]~25 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][6]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_21_add_1_o[6]~24 ),
	.combout(\u1_m0_wo0_mtree_mult1_21_add_1_o[7]~25_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_21_add_1_o[7]~26 ));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[7]~25 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[7]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_21_add_1_o[8]~27 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][8]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_21_add_1_o[7]~26 ),
	.combout(\u1_m0_wo0_mtree_mult1_21_add_1_o[8]~27_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_21_add_1_o[8]~28 ));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[8]~27 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[8]~27 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_21_add_1_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_21_add_1_o[8]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_21_add_1_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_2_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_2_o[8]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_2_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_21_add_1_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_21_add_1_o[7]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_21_add_1_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_2_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_2_o[7]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_2_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_21_add_1_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_21_add_1_o[6]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_21_add_1_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_2_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_2_o[6]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_2_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_21_add_1_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_21_add_1_o[5]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_21_add_1_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_2_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_2_o[5]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_2_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_21_add_1_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_21_add_1_o[4]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_21_add_1_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_2_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_2_o[4]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_2_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_21_add_1_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_21_add_1_o[3]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_21_add_1_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_2_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_2_o[3]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_2_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_21_add_1_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_21_add_1_o[2]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_21_add_1_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_2_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_2_o[2]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_2_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_21_add_1_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_21_add_1_o[1]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_21_add_1_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_0_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_0_o[1]~12_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_0_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_2_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_0_o[1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_2_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_21_add_1_o[0] (
	.clk(clk),
	.d(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_21_add_1_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_10_o[1]~15 (
	.dataa(\u1_m0_wo0_mtree_mult1_20_sub_2_o[1]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_21_add_1_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_add0_10_o[1]~15_combout ),
	.cout(\u1_m0_wo0_mtree_add0_10_o[1]~16 ));
defparam \u1_m0_wo0_mtree_add0_10_o[1]~15 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_add0_10_o[1]~15 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_10_o[2]~17 (
	.dataa(\u1_m0_wo0_mtree_mult1_20_sub_2_o[2]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_21_add_1_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_10_o[1]~16 ),
	.combout(\u1_m0_wo0_mtree_add0_10_o[2]~17_combout ),
	.cout(\u1_m0_wo0_mtree_add0_10_o[2]~18 ));
defparam \u1_m0_wo0_mtree_add0_10_o[2]~17 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_10_o[2]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_10_o[3]~19 (
	.dataa(\u1_m0_wo0_mtree_mult1_20_sub_2_o[3]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_21_add_1_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_10_o[2]~18 ),
	.combout(\u1_m0_wo0_mtree_add0_10_o[3]~19_combout ),
	.cout(\u1_m0_wo0_mtree_add0_10_o[3]~20 ));
defparam \u1_m0_wo0_mtree_add0_10_o[3]~19 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_10_o[3]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_10_o[4]~21 (
	.dataa(\u1_m0_wo0_mtree_mult1_20_sub_2_o[4]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_21_add_1_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_10_o[3]~20 ),
	.combout(\u1_m0_wo0_mtree_add0_10_o[4]~21_combout ),
	.cout(\u1_m0_wo0_mtree_add0_10_o[4]~22 ));
defparam \u1_m0_wo0_mtree_add0_10_o[4]~21 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_10_o[4]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_10_o[5]~23 (
	.dataa(\u1_m0_wo0_mtree_mult1_20_sub_2_o[5]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_21_add_1_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_10_o[4]~22 ),
	.combout(\u1_m0_wo0_mtree_add0_10_o[5]~23_combout ),
	.cout(\u1_m0_wo0_mtree_add0_10_o[5]~24 ));
defparam \u1_m0_wo0_mtree_add0_10_o[5]~23 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_10_o[5]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_10_o[6]~25 (
	.dataa(\u1_m0_wo0_mtree_mult1_20_sub_2_o[6]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_21_add_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_10_o[5]~24 ),
	.combout(\u1_m0_wo0_mtree_add0_10_o[6]~25_combout ),
	.cout(\u1_m0_wo0_mtree_add0_10_o[6]~26 ));
defparam \u1_m0_wo0_mtree_add0_10_o[6]~25 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_10_o[6]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_10_o[7]~27 (
	.dataa(\u1_m0_wo0_mtree_mult1_20_sub_2_o[7]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_21_add_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_10_o[6]~26 ),
	.combout(\u1_m0_wo0_mtree_add0_10_o[7]~27_combout ),
	.cout(\u1_m0_wo0_mtree_add0_10_o[7]~28 ));
defparam \u1_m0_wo0_mtree_add0_10_o[7]~27 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_10_o[7]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_10_o[8]~29 (
	.dataa(\u1_m0_wo0_mtree_mult1_20_sub_2_o[8]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_21_add_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_10_o[7]~28 ),
	.combout(\u1_m0_wo0_mtree_add0_10_o[8]~29_combout ),
	.cout(\u1_m0_wo0_mtree_add0_10_o[8]~30 ));
defparam \u1_m0_wo0_mtree_add0_10_o[8]~29 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_10_o[8]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_10_o[9]~31 (
	.dataa(\u1_m0_wo0_mtree_mult1_20_sub_2_o[9]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_21_add_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_10_o[8]~30 ),
	.combout(\u1_m0_wo0_mtree_add0_10_o[9]~31_combout ),
	.cout(\u1_m0_wo0_mtree_add0_10_o[9]~32 ));
defparam \u1_m0_wo0_mtree_add0_10_o[9]~31 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_10_o[9]~31 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add0_10_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_10_o[9]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_10_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_10_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_10_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_22_sub_1_o[2]~13 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][0]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[2]~13_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[2]~14 ));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[2]~13 .lut_mask = 16'h66DD;
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[2]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_22_sub_1_o[3]~15 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][1]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_22_sub_1_o[2]~14 ),
	.combout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[3]~15_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[3]~16 ));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[3]~15 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[3]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_22_sub_1_o[4]~17 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][2]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_22_sub_1_o[3]~16 ),
	.combout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[4]~17_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[4]~18 ));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[4]~17 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[4]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_22_sub_1_o[5]~19 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][3]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_22_sub_1_o[4]~18 ),
	.combout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[5]~19_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[5]~20 ));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[5]~19 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[5]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_22_sub_1_o[6]~21 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][4]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_22_sub_1_o[5]~20 ),
	.combout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[6]~21_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[6]~22 ));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[6]~21 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[6]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_22_sub_1_o[7]~23 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][5]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_22_sub_1_o[6]~22 ),
	.combout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[7]~23_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[7]~24 ));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[7]~23 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[7]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_22_sub_1_o[8]~25 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][6]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_22_sub_1_o[7]~24 ),
	.combout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[8]~25_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[8]~26 ));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[8]~25 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[8]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_22_sub_1_o[9]~27 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][7]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_22_sub_1_o[8]~26 ),
	.combout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[9]~27_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[9]~28 ));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[9]~27 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[9]~27 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_22_sub_1_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_22_sub_1_o[9]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_22_sub_1_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_10_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_10_o[8]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_10_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_10_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_10_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_22_sub_1_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_22_sub_1_o[8]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_22_sub_1_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_10_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_10_o[7]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_10_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_10_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_10_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_22_sub_1_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_22_sub_1_o[7]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_22_sub_1_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_10_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_10_o[6]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_10_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_10_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_10_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_22_sub_1_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_22_sub_1_o[6]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_22_sub_1_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_10_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_10_o[5]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_10_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_10_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_10_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_22_sub_1_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_22_sub_1_o[5]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_22_sub_1_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_10_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_10_o[4]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_10_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_10_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_10_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_22_sub_1_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_22_sub_1_o[4]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_22_sub_1_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_10_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_10_o[3]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_10_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_10_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_10_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_22_sub_1_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_22_sub_1_o[3]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_22_sub_1_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_10_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_10_o[2]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_10_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_10_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_10_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_22_sub_1_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_22_sub_1_o[2]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_22_sub_1_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_10_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_10_o[1]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_10_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_10_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_10_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_22_sub_1_o[1] (
	.clk(clk),
	.d(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_22_sub_1_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_2_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_0_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_2_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_10_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_2_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_10_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_10_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_10_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_22_sub_1_o[0] (
	.clk(clk),
	.d(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_22_sub_1_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_5_o[0]~17 (
	.dataa(\u1_m0_wo0_mtree_add0_10_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_22_sub_1_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_add1_5_o[0]~17_combout ),
	.cout(\u1_m0_wo0_mtree_add1_5_o[0]~18 ));
defparam \u1_m0_wo0_mtree_add1_5_o[0]~17 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_add1_5_o[0]~17 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_5_o[1]~19 (
	.dataa(\u1_m0_wo0_mtree_add0_10_o[1]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_22_sub_1_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_5_o[0]~18 ),
	.combout(\u1_m0_wo0_mtree_add1_5_o[1]~19_combout ),
	.cout(\u1_m0_wo0_mtree_add1_5_o[1]~20 ));
defparam \u1_m0_wo0_mtree_add1_5_o[1]~19 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_5_o[1]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_5_o[2]~21 (
	.dataa(\u1_m0_wo0_mtree_add0_10_o[2]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_22_sub_1_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_5_o[1]~20 ),
	.combout(\u1_m0_wo0_mtree_add1_5_o[2]~21_combout ),
	.cout(\u1_m0_wo0_mtree_add1_5_o[2]~22 ));
defparam \u1_m0_wo0_mtree_add1_5_o[2]~21 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_5_o[2]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_5_o[3]~23 (
	.dataa(\u1_m0_wo0_mtree_add0_10_o[3]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_22_sub_1_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_5_o[2]~22 ),
	.combout(\u1_m0_wo0_mtree_add1_5_o[3]~23_combout ),
	.cout(\u1_m0_wo0_mtree_add1_5_o[3]~24 ));
defparam \u1_m0_wo0_mtree_add1_5_o[3]~23 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_5_o[3]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_5_o[4]~25 (
	.dataa(\u1_m0_wo0_mtree_add0_10_o[4]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_22_sub_1_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_5_o[3]~24 ),
	.combout(\u1_m0_wo0_mtree_add1_5_o[4]~25_combout ),
	.cout(\u1_m0_wo0_mtree_add1_5_o[4]~26 ));
defparam \u1_m0_wo0_mtree_add1_5_o[4]~25 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_5_o[4]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_5_o[5]~27 (
	.dataa(\u1_m0_wo0_mtree_add0_10_o[5]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_22_sub_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_5_o[4]~26 ),
	.combout(\u1_m0_wo0_mtree_add1_5_o[5]~27_combout ),
	.cout(\u1_m0_wo0_mtree_add1_5_o[5]~28 ));
defparam \u1_m0_wo0_mtree_add1_5_o[5]~27 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_5_o[5]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_5_o[6]~29 (
	.dataa(\u1_m0_wo0_mtree_add0_10_o[6]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_22_sub_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_5_o[5]~28 ),
	.combout(\u1_m0_wo0_mtree_add1_5_o[6]~29_combout ),
	.cout(\u1_m0_wo0_mtree_add1_5_o[6]~30 ));
defparam \u1_m0_wo0_mtree_add1_5_o[6]~29 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_5_o[6]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_5_o[7]~31 (
	.dataa(\u1_m0_wo0_mtree_add0_10_o[7]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_22_sub_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_5_o[6]~30 ),
	.combout(\u1_m0_wo0_mtree_add1_5_o[7]~31_combout ),
	.cout(\u1_m0_wo0_mtree_add1_5_o[7]~32 ));
defparam \u1_m0_wo0_mtree_add1_5_o[7]~31 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_5_o[7]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_5_o[8]~33 (
	.dataa(\u1_m0_wo0_mtree_add0_10_o[8]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_22_sub_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_5_o[7]~32 ),
	.combout(\u1_m0_wo0_mtree_add1_5_o[8]~33_combout ),
	.cout(\u1_m0_wo0_mtree_add1_5_o[8]~34 ));
defparam \u1_m0_wo0_mtree_add1_5_o[8]~33 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_5_o[8]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_5_o[9]~35 (
	.dataa(\u1_m0_wo0_mtree_add0_10_o[9]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_22_sub_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_5_o[8]~34 ),
	.combout(\u1_m0_wo0_mtree_add1_5_o[9]~35_combout ),
	.cout(\u1_m0_wo0_mtree_add1_5_o[9]~36 ));
defparam \u1_m0_wo0_mtree_add1_5_o[9]~35 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_5_o[9]~35 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add1_5_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_5_o[9]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_5_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_5_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_5_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_4_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[8]~36_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_5_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_5_o[8]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_5_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_5_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_5_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_4_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[7]~34_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_5_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_5_o[7]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_5_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_5_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_5_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_4_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[6]~32_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_5_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_5_o[6]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_5_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_5_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_5_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_4_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[5]~30_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_5_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_5_o[5]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_5_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_5_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_5_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_4_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[4]~28_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_5_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_5_o[4]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_5_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_5_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_5_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_4_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[3]~26_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_5_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_5_o[3]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_5_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_5_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_5_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_4_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[2]~24_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_5_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_5_o[2]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_5_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_5_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_5_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_4_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[1]~22_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_5_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_5_o[1]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_5_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_5_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_5_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_4_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[0]~20_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_5_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_5_o[0]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_5_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_5_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_5_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[0]~21 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_add2_2_o[0]~21_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[0]~22 ));
defparam \u1_m0_wo0_mtree_add2_2_o[0]~21 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_add2_2_o[0]~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[1]~23 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[1]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_2_o[0]~22 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[1]~23_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[1]~24 ));
defparam \u1_m0_wo0_mtree_add2_2_o[1]~23 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_2_o[1]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[2]~25 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[2]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_2_o[1]~24 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[2]~25_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[2]~26 ));
defparam \u1_m0_wo0_mtree_add2_2_o[2]~25 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add2_2_o[2]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[3]~27 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[3]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_2_o[2]~26 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[3]~27_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[3]~28 ));
defparam \u1_m0_wo0_mtree_add2_2_o[3]~27 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_2_o[3]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[4]~29 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[4]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_2_o[3]~28 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[4]~29_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[4]~30 ));
defparam \u1_m0_wo0_mtree_add2_2_o[4]~29 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add2_2_o[4]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[5]~31 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[5]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_2_o[4]~30 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[5]~31_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[5]~32 ));
defparam \u1_m0_wo0_mtree_add2_2_o[5]~31 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_2_o[5]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[6]~33 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[6]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_2_o[5]~32 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[6]~33_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[6]~34 ));
defparam \u1_m0_wo0_mtree_add2_2_o[6]~33 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add2_2_o[6]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[7]~35 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[7]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_2_o[6]~34 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[7]~35_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[7]~36 ));
defparam \u1_m0_wo0_mtree_add2_2_o[7]~35 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_2_o[7]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[8]~37 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[8]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_2_o[7]~36 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[8]~37_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[8]~38 ));
defparam \u1_m0_wo0_mtree_add2_2_o[8]~37 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add2_2_o[8]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[9]~39 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[9]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_2_o[8]~38 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[9]~39_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[9]~40 ));
defparam \u1_m0_wo0_mtree_add2_2_o[9]~39 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_2_o[9]~39 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add2_2_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[9]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_25_sub_0_o[1]~12 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][0]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[1]~12_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[1]~13 ));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[1]~12 .lut_mask = 16'h6611;
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[1]~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_25_sub_0_o[2]~14 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_25_sub_0_o[1]~13 ),
	.combout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[2]~14_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[2]~15 ));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[2]~14 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[2]~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_25_sub_0_o[3]~16 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_25_sub_0_o[2]~15 ),
	.combout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[3]~16_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[3]~17 ));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[3]~16 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[3]~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_25_sub_0_o[4]~18 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_25_sub_0_o[3]~17 ),
	.combout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[4]~18_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[4]~19 ));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[4]~18 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[4]~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_25_sub_0_o[5]~20 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_25_sub_0_o[4]~19 ),
	.combout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[5]~20_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[5]~21 ));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[5]~20 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[5]~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_25_sub_0_o[6]~22 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_25_sub_0_o[5]~21 ),
	.combout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[6]~22_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[6]~23 ));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[6]~22 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[6]~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_25_sub_0_o[7]~24 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_25_sub_0_o[6]~23 ),
	.combout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[7]~24_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[7]~25 ));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[7]~24 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[7]~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_25_sub_0_o[8]~26 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_25_sub_0_o[7]~25 ),
	.combout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[8]~26_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[8]~27 ));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[8]~26 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[8]~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_25_sub_0_o[9]~28 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_25_sub_0_o[8]~27 ),
	.combout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[9]~28_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[9]~29 ));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[9]~28 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[9]~28 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_25_sub_0_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_25_sub_0_o[9]~28_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_25_sub_0_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_25_sub_0_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_25_sub_0_o[8]~26_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_25_sub_0_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_25_sub_0_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_25_sub_0_o[7]~24_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_25_sub_0_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_25_sub_0_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_25_sub_0_o[6]~22_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_25_sub_0_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_25_sub_0_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_25_sub_0_o[5]~20_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_25_sub_0_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_25_sub_0_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_25_sub_0_o[4]~18_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_25_sub_0_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_25_sub_0_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_25_sub_0_o[3]~16_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_25_sub_0_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_25_sub_0_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_25_sub_0_o[2]~14_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_25_sub_0_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_25_sub_0_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_25_sub_0_o[1]~12_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_25_sub_0_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_25_sub_0_o[0] (
	.clk(clk),
	.d(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_25_sub_0_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_12_o[0]~14 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][0]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_25_sub_0_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_add0_12_o[0]~14_combout ),
	.cout(\u1_m0_wo0_mtree_add0_12_o[0]~15 ));
defparam \u1_m0_wo0_mtree_add0_12_o[0]~14 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_add0_12_o[0]~14 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_12_o[1]~16 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][1]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_25_sub_0_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_12_o[0]~15 ),
	.combout(\u1_m0_wo0_mtree_add0_12_o[1]~16_combout ),
	.cout(\u1_m0_wo0_mtree_add0_12_o[1]~17 ));
defparam \u1_m0_wo0_mtree_add0_12_o[1]~16 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_12_o[1]~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_12_o[2]~18 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][2]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_25_sub_0_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_12_o[1]~17 ),
	.combout(\u1_m0_wo0_mtree_add0_12_o[2]~18_combout ),
	.cout(\u1_m0_wo0_mtree_add0_12_o[2]~19 ));
defparam \u1_m0_wo0_mtree_add0_12_o[2]~18 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_12_o[2]~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_12_o[3]~20 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][3]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_25_sub_0_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_12_o[2]~19 ),
	.combout(\u1_m0_wo0_mtree_add0_12_o[3]~20_combout ),
	.cout(\u1_m0_wo0_mtree_add0_12_o[3]~21 ));
defparam \u1_m0_wo0_mtree_add0_12_o[3]~20 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_12_o[3]~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_12_o[4]~22 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][4]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_25_sub_0_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_12_o[3]~21 ),
	.combout(\u1_m0_wo0_mtree_add0_12_o[4]~22_combout ),
	.cout(\u1_m0_wo0_mtree_add0_12_o[4]~23 ));
defparam \u1_m0_wo0_mtree_add0_12_o[4]~22 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_12_o[4]~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_12_o[5]~24 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][5]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_25_sub_0_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_12_o[4]~23 ),
	.combout(\u1_m0_wo0_mtree_add0_12_o[5]~24_combout ),
	.cout(\u1_m0_wo0_mtree_add0_12_o[5]~25 ));
defparam \u1_m0_wo0_mtree_add0_12_o[5]~24 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_12_o[5]~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_12_o[6]~26 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][6]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_25_sub_0_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_12_o[5]~25 ),
	.combout(\u1_m0_wo0_mtree_add0_12_o[6]~26_combout ),
	.cout(\u1_m0_wo0_mtree_add0_12_o[6]~27 ));
defparam \u1_m0_wo0_mtree_add0_12_o[6]~26 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_12_o[6]~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_12_o[7]~28 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][7]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_25_sub_0_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_12_o[6]~27 ),
	.combout(\u1_m0_wo0_mtree_add0_12_o[7]~28_combout ),
	.cout(\u1_m0_wo0_mtree_add0_12_o[7]~29 ));
defparam \u1_m0_wo0_mtree_add0_12_o[7]~28 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_12_o[7]~28 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_12_o[8]~30 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][8]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_25_sub_0_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_12_o[7]~29 ),
	.combout(\u1_m0_wo0_mtree_add0_12_o[8]~30_combout ),
	.cout(\u1_m0_wo0_mtree_add0_12_o[8]~31 ));
defparam \u1_m0_wo0_mtree_add0_12_o[8]~30 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_12_o[8]~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_12_o[9]~32 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][9]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_25_sub_0_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_12_o[8]~31 ),
	.combout(\u1_m0_wo0_mtree_add0_12_o[9]~32_combout ),
	.cout(\u1_m0_wo0_mtree_add0_12_o[9]~33 ));
defparam \u1_m0_wo0_mtree_add0_12_o[9]~32 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_12_o[9]~32 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add0_12_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_12_o[9]~32_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_12_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_12_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_12_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_2_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[8]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_12_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_12_o[8]~30_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_12_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_12_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_12_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_2_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[7]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_12_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_12_o[7]~28_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_12_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_12_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_12_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_2_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[6]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_12_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_12_o[6]~26_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_12_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_12_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_12_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_2_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[5]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_12_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_12_o[5]~24_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_12_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_12_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_12_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_2_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[4]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_12_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_12_o[4]~22_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_12_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_12_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_12_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_2_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[3]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_12_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_12_o[3]~20_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_12_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_12_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_12_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_2_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[2]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_12_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_12_o[2]~18_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_12_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_12_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_12_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_2_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[1]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_12_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_12_o[1]~16_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_12_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_12_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_12_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_2_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[0]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_12_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_12_o[0]~14_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_12_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_12_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_12_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[0]~21 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u1_m0_wo0_mtree_add3_1_o[0]~21_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[0]~22 ));
defparam \u1_m0_wo0_mtree_add3_1_o[0]~21 .lut_mask = 16'h6688;
defparam \u1_m0_wo0_mtree_add3_1_o[0]~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[1]~23 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[1]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_1_o[0]~22 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[1]~23_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[1]~24 ));
defparam \u1_m0_wo0_mtree_add3_1_o[1]~23 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_1_o[1]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[2]~25 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[2]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_1_o[1]~24 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[2]~25_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[2]~26 ));
defparam \u1_m0_wo0_mtree_add3_1_o[2]~25 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add3_1_o[2]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[3]~27 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[3]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_1_o[2]~26 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[3]~27_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[3]~28 ));
defparam \u1_m0_wo0_mtree_add3_1_o[3]~27 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_1_o[3]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[4]~29 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[4]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_1_o[3]~28 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[4]~29_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[4]~30 ));
defparam \u1_m0_wo0_mtree_add3_1_o[4]~29 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add3_1_o[4]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[5]~31 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[5]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_1_o[4]~30 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[5]~31_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[5]~32 ));
defparam \u1_m0_wo0_mtree_add3_1_o[5]~31 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_1_o[5]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[6]~33 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[6]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_1_o[5]~32 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[6]~33_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[6]~34 ));
defparam \u1_m0_wo0_mtree_add3_1_o[6]~33 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add3_1_o[6]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[7]~35 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[7]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_1_o[6]~34 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[7]~35_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[7]~36 ));
defparam \u1_m0_wo0_mtree_add3_1_o[7]~35 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_1_o[7]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[8]~37 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[8]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_1_o[7]~36 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[8]~37_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[8]~38 ));
defparam \u1_m0_wo0_mtree_add3_1_o[8]~37 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add3_1_o[8]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[9]~39 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[9]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_1_o[8]~38 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[9]~39_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[9]~40 ));
defparam \u1_m0_wo0_mtree_add3_1_o[9]~39 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_1_o[9]~39 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add3_1_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[9]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[9] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_0_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[8]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_1_o[8] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[8]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[8]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[8] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[8] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_0_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[7]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_1_o[7] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[7]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[7]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[7] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[7] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_0_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[6]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_1_o[6] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[6]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[6]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[6] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[6] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_0_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[5]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_1_o[5] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[5]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[5]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[5] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[5] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_0_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[4]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_1_o[4] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[4]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[4]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[4] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[4] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_0_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[3]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_1_o[3] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[3]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[3]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[3] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[3] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_0_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[2]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_1_o[2] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[2]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[2]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[2] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[2] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_0_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[1]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_1_o[1] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[1]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[1]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[1] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[1] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_0_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[0]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[0] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_1_o[0] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[0]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[0]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[0] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[9]~13 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[0]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\u1_m0_wo0_mtree_add4_0_o[9]~13_cout ));
defparam \u1_m0_wo0_mtree_add4_0_o[9]~13 .lut_mask = 16'h0088;
defparam \u1_m0_wo0_mtree_add4_0_o[9]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[9]~15 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[1]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add4_0_o[9]~13_cout ),
	.combout(),
	.cout(\u1_m0_wo0_mtree_add4_0_o[9]~15_cout ));
defparam \u1_m0_wo0_mtree_add4_0_o[9]~15 .lut_mask = 16'h0017;
defparam \u1_m0_wo0_mtree_add4_0_o[9]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[9]~17 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[2]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add4_0_o[9]~15_cout ),
	.combout(),
	.cout(\u1_m0_wo0_mtree_add4_0_o[9]~17_cout ));
defparam \u1_m0_wo0_mtree_add4_0_o[9]~17 .lut_mask = 16'h008E;
defparam \u1_m0_wo0_mtree_add4_0_o[9]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[9]~19 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[3]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add4_0_o[9]~17_cout ),
	.combout(),
	.cout(\u1_m0_wo0_mtree_add4_0_o[9]~19_cout ));
defparam \u1_m0_wo0_mtree_add4_0_o[9]~19 .lut_mask = 16'h0017;
defparam \u1_m0_wo0_mtree_add4_0_o[9]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[9]~21 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[4]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add4_0_o[9]~19_cout ),
	.combout(),
	.cout(\u1_m0_wo0_mtree_add4_0_o[9]~21_cout ));
defparam \u1_m0_wo0_mtree_add4_0_o[9]~21 .lut_mask = 16'h008E;
defparam \u1_m0_wo0_mtree_add4_0_o[9]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[9]~23 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[5]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add4_0_o[9]~21_cout ),
	.combout(),
	.cout(\u1_m0_wo0_mtree_add4_0_o[9]~23_cout ));
defparam \u1_m0_wo0_mtree_add4_0_o[9]~23 .lut_mask = 16'h0017;
defparam \u1_m0_wo0_mtree_add4_0_o[9]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[9]~25 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[6]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add4_0_o[9]~23_cout ),
	.combout(),
	.cout(\u1_m0_wo0_mtree_add4_0_o[9]~25_cout ));
defparam \u1_m0_wo0_mtree_add4_0_o[9]~25 .lut_mask = 16'h008E;
defparam \u1_m0_wo0_mtree_add4_0_o[9]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[9]~27 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[7]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add4_0_o[9]~25_cout ),
	.combout(),
	.cout(\u1_m0_wo0_mtree_add4_0_o[9]~27_cout ));
defparam \u1_m0_wo0_mtree_add4_0_o[9]~27 .lut_mask = 16'h0017;
defparam \u1_m0_wo0_mtree_add4_0_o[9]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[9]~29 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[8]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add4_0_o[9]~27_cout ),
	.combout(),
	.cout(\u1_m0_wo0_mtree_add4_0_o[9]~29_cout ));
defparam \u1_m0_wo0_mtree_add4_0_o[9]~29 .lut_mask = 16'h008E;
defparam \u1_m0_wo0_mtree_add4_0_o[9]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[9]~30 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[9]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add4_0_o[9]~29_cout ),
	.combout(\u1_m0_wo0_mtree_add4_0_o[9]~30_combout ),
	.cout(\u1_m0_wo0_mtree_add4_0_o[9]~31 ));
defparam \u1_m0_wo0_mtree_add4_0_o[9]~30 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add4_0_o[9]~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_5_sub_0_o[1]~12 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][0]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[1]~12_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[1]~13 ));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[1]~12 .lut_mask = 16'h6611;
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[1]~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_5_sub_0_o[2]~14 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_5_sub_0_o[1]~13 ),
	.combout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[2]~14_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[2]~15 ));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[2]~14 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[2]~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_5_sub_0_o[3]~16 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_5_sub_0_o[2]~15 ),
	.combout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[3]~16_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[3]~17 ));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[3]~16 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[3]~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_5_sub_0_o[4]~18 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_5_sub_0_o[3]~17 ),
	.combout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[4]~18_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[4]~19 ));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[4]~18 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[4]~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_5_sub_0_o[5]~20 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_5_sub_0_o[4]~19 ),
	.combout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[5]~20_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[5]~21 ));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[5]~20 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[5]~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_5_sub_0_o[6]~22 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_5_sub_0_o[5]~21 ),
	.combout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[6]~22_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[6]~23 ));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[6]~22 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[6]~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_5_sub_0_o[7]~24 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_5_sub_0_o[6]~23 ),
	.combout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[7]~24_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[7]~25 ));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[7]~24 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[7]~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_5_sub_0_o[8]~26 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_5_sub_0_o[7]~25 ),
	.combout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[8]~26_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[8]~27 ));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[8]~26 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[8]~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_5_sub_0_o[9]~28 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_5_sub_0_o[8]~27 ),
	.combout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[9]~28_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[9]~29 ));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[9]~28 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[9]~28 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_5_sub_0_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_5_sub_0_o[9]~28_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_5_sub_0_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_5_sub_0_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_5_sub_0_o[8]~26_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_5_sub_0_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_5_sub_0_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_5_sub_0_o[7]~24_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_5_sub_0_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_5_sub_0_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_5_sub_0_o[6]~22_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_5_sub_0_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_5_sub_0_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_5_sub_0_o[5]~20_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_5_sub_0_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_5_sub_0_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_5_sub_0_o[4]~18_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_5_sub_0_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_5_sub_0_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_5_sub_0_o[3]~16_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_5_sub_0_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_5_sub_0_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_5_sub_0_o[2]~14_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_5_sub_0_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_5_sub_0_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_5_sub_0_o[1]~12_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_5_sub_0_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_5_sub_0_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_5_sub_0_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_1_o[0]~14 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][0]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_5_sub_0_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_add1_1_o[0]~14_combout ),
	.cout(\u0_m0_wo0_mtree_add1_1_o[0]~15 ));
defparam \u0_m0_wo0_mtree_add1_1_o[0]~14 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_add1_1_o[0]~14 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_1_o[1]~16 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][1]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_5_sub_0_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_1_o[0]~15 ),
	.combout(\u0_m0_wo0_mtree_add1_1_o[1]~16_combout ),
	.cout(\u0_m0_wo0_mtree_add1_1_o[1]~17 ));
defparam \u0_m0_wo0_mtree_add1_1_o[1]~16 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_1_o[1]~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_1_o[2]~18 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][2]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_5_sub_0_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_1_o[1]~17 ),
	.combout(\u0_m0_wo0_mtree_add1_1_o[2]~18_combout ),
	.cout(\u0_m0_wo0_mtree_add1_1_o[2]~19 ));
defparam \u0_m0_wo0_mtree_add1_1_o[2]~18 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_1_o[2]~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_1_o[3]~20 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][3]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_5_sub_0_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_1_o[2]~19 ),
	.combout(\u0_m0_wo0_mtree_add1_1_o[3]~20_combout ),
	.cout(\u0_m0_wo0_mtree_add1_1_o[3]~21 ));
defparam \u0_m0_wo0_mtree_add1_1_o[3]~20 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_1_o[3]~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_1_o[4]~22 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][4]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_5_sub_0_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_1_o[3]~21 ),
	.combout(\u0_m0_wo0_mtree_add1_1_o[4]~22_combout ),
	.cout(\u0_m0_wo0_mtree_add1_1_o[4]~23 ));
defparam \u0_m0_wo0_mtree_add1_1_o[4]~22 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_1_o[4]~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_1_o[5]~24 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][5]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_5_sub_0_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_1_o[4]~23 ),
	.combout(\u0_m0_wo0_mtree_add1_1_o[5]~24_combout ),
	.cout(\u0_m0_wo0_mtree_add1_1_o[5]~25 ));
defparam \u0_m0_wo0_mtree_add1_1_o[5]~24 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_1_o[5]~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_1_o[6]~26 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][6]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_5_sub_0_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_1_o[5]~25 ),
	.combout(\u0_m0_wo0_mtree_add1_1_o[6]~26_combout ),
	.cout(\u0_m0_wo0_mtree_add1_1_o[6]~27 ));
defparam \u0_m0_wo0_mtree_add1_1_o[6]~26 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_1_o[6]~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_1_o[7]~28 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][7]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_5_sub_0_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_1_o[6]~27 ),
	.combout(\u0_m0_wo0_mtree_add1_1_o[7]~28_combout ),
	.cout(\u0_m0_wo0_mtree_add1_1_o[7]~29 ));
defparam \u0_m0_wo0_mtree_add1_1_o[7]~28 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_1_o[7]~28 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_1_o[8]~30 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][8]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_5_sub_0_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_1_o[7]~29 ),
	.combout(\u0_m0_wo0_mtree_add1_1_o[8]~30_combout ),
	.cout(\u0_m0_wo0_mtree_add1_1_o[8]~31 ));
defparam \u0_m0_wo0_mtree_add1_1_o[8]~30 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_1_o[8]~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_1_o[9]~32 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][9]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_5_sub_0_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_1_o[8]~31 ),
	.combout(\u0_m0_wo0_mtree_add1_1_o[9]~32_combout ),
	.cout(\u0_m0_wo0_mtree_add1_1_o[9]~33 ));
defparam \u0_m0_wo0_mtree_add1_1_o[9]~32 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_1_o[9]~32 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add1_1_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_1_o[9]~32_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_1_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_1_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_1_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_8_sub_1_o[2]~13 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][0]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[2]~13_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[2]~14 ));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[2]~13 .lut_mask = 16'h66DD;
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[2]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_8_sub_1_o[3]~15 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][1]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_8_sub_1_o[2]~14 ),
	.combout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[3]~15_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[3]~16 ));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[3]~15 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[3]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_8_sub_1_o[4]~17 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][2]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_8_sub_1_o[3]~16 ),
	.combout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[4]~17_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[4]~18 ));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[4]~17 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[4]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_8_sub_1_o[5]~19 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][3]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_8_sub_1_o[4]~18 ),
	.combout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[5]~19_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[5]~20 ));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[5]~19 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[5]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_8_sub_1_o[6]~21 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][4]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_8_sub_1_o[5]~20 ),
	.combout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[6]~21_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[6]~22 ));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[6]~21 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[6]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_8_sub_1_o[7]~23 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][5]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_8_sub_1_o[6]~22 ),
	.combout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[7]~23_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[7]~24 ));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[7]~23 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[7]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_8_sub_1_o[8]~25 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][6]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_8_sub_1_o[7]~24 ),
	.combout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[8]~25_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[8]~26 ));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[8]~25 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[8]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_8_sub_1_o[9]~27 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][7]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_8_sub_1_o[8]~26 ),
	.combout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[9]~27_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[9]~28 ));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[9]~27 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[9]~27 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_8_sub_1_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_8_sub_1_o[9]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_8_sub_1_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_9_add_1_o[1]~13 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][0]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_9_add_1_o[1]~13_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_9_add_1_o[1]~14 ));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[1]~13 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[1]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_9_add_1_o[2]~15 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][2]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_9_add_1_o[1]~14 ),
	.combout(\u0_m0_wo0_mtree_mult1_9_add_1_o[2]~15_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_9_add_1_o[2]~16 ));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[2]~15 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[2]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_9_add_1_o[3]~17 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][2]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_9_add_1_o[2]~16 ),
	.combout(\u0_m0_wo0_mtree_mult1_9_add_1_o[3]~17_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_9_add_1_o[3]~18 ));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[3]~17 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[3]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_9_add_1_o[4]~19 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][4]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_9_add_1_o[3]~18 ),
	.combout(\u0_m0_wo0_mtree_mult1_9_add_1_o[4]~19_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_9_add_1_o[4]~20 ));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[4]~19 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[4]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_9_add_1_o[5]~21 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][4]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_9_add_1_o[4]~20 ),
	.combout(\u0_m0_wo0_mtree_mult1_9_add_1_o[5]~21_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_9_add_1_o[5]~22 ));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[5]~21 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[5]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_9_add_1_o[6]~23 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][6]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_9_add_1_o[5]~22 ),
	.combout(\u0_m0_wo0_mtree_mult1_9_add_1_o[6]~23_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_9_add_1_o[6]~24 ));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[6]~23 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[6]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_9_add_1_o[7]~25 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][6]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_9_add_1_o[6]~24 ),
	.combout(\u0_m0_wo0_mtree_mult1_9_add_1_o[7]~25_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_9_add_1_o[7]~26 ));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[7]~25 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[7]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_9_add_1_o[8]~27 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][8]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_9_add_1_o[7]~26 ),
	.combout(\u0_m0_wo0_mtree_mult1_9_add_1_o[8]~27_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_9_add_1_o[8]~28 ));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[8]~27 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[8]~27 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_9_add_1_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_9_add_1_o[8]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_9_add_1_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_8_sub_1_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_8_sub_1_o[8]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_8_sub_1_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_9_add_1_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_9_add_1_o[7]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_9_add_1_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_8_sub_1_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_8_sub_1_o[7]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_8_sub_1_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_9_add_1_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_9_add_1_o[6]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_9_add_1_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_8_sub_1_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_8_sub_1_o[6]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_8_sub_1_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_9_add_1_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_9_add_1_o[5]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_9_add_1_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_8_sub_1_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_8_sub_1_o[5]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_8_sub_1_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_9_add_1_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_9_add_1_o[4]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_9_add_1_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_8_sub_1_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_8_sub_1_o[4]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_8_sub_1_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_9_add_1_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_9_add_1_o[3]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_9_add_1_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_8_sub_1_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_8_sub_1_o[3]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_8_sub_1_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_9_add_1_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_9_add_1_o[2]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_9_add_1_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_8_sub_1_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_8_sub_1_o[2]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_8_sub_1_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_9_add_1_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_9_add_1_o[1]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_9_add_1_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_8_sub_1_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_8_sub_1_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_9_add_1_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_9_add_1_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_4_o[1]~15 (
	.dataa(\u0_m0_wo0_mtree_mult1_8_sub_1_o[1]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_9_add_1_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_add0_4_o[1]~15_combout ),
	.cout(\u0_m0_wo0_mtree_add0_4_o[1]~16 ));
defparam \u0_m0_wo0_mtree_add0_4_o[1]~15 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_add0_4_o[1]~15 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_4_o[2]~17 (
	.dataa(\u0_m0_wo0_mtree_mult1_8_sub_1_o[2]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_9_add_1_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_4_o[1]~16 ),
	.combout(\u0_m0_wo0_mtree_add0_4_o[2]~17_combout ),
	.cout(\u0_m0_wo0_mtree_add0_4_o[2]~18 ));
defparam \u0_m0_wo0_mtree_add0_4_o[2]~17 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_4_o[2]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_4_o[3]~19 (
	.dataa(\u0_m0_wo0_mtree_mult1_8_sub_1_o[3]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_9_add_1_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_4_o[2]~18 ),
	.combout(\u0_m0_wo0_mtree_add0_4_o[3]~19_combout ),
	.cout(\u0_m0_wo0_mtree_add0_4_o[3]~20 ));
defparam \u0_m0_wo0_mtree_add0_4_o[3]~19 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_4_o[3]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_4_o[4]~21 (
	.dataa(\u0_m0_wo0_mtree_mult1_8_sub_1_o[4]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_9_add_1_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_4_o[3]~20 ),
	.combout(\u0_m0_wo0_mtree_add0_4_o[4]~21_combout ),
	.cout(\u0_m0_wo0_mtree_add0_4_o[4]~22 ));
defparam \u0_m0_wo0_mtree_add0_4_o[4]~21 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_4_o[4]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_4_o[5]~23 (
	.dataa(\u0_m0_wo0_mtree_mult1_8_sub_1_o[5]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_9_add_1_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_4_o[4]~22 ),
	.combout(\u0_m0_wo0_mtree_add0_4_o[5]~23_combout ),
	.cout(\u0_m0_wo0_mtree_add0_4_o[5]~24 ));
defparam \u0_m0_wo0_mtree_add0_4_o[5]~23 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_4_o[5]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_4_o[6]~25 (
	.dataa(\u0_m0_wo0_mtree_mult1_8_sub_1_o[6]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_9_add_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_4_o[5]~24 ),
	.combout(\u0_m0_wo0_mtree_add0_4_o[6]~25_combout ),
	.cout(\u0_m0_wo0_mtree_add0_4_o[6]~26 ));
defparam \u0_m0_wo0_mtree_add0_4_o[6]~25 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_4_o[6]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_4_o[7]~27 (
	.dataa(\u0_m0_wo0_mtree_mult1_8_sub_1_o[7]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_9_add_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_4_o[6]~26 ),
	.combout(\u0_m0_wo0_mtree_add0_4_o[7]~27_combout ),
	.cout(\u0_m0_wo0_mtree_add0_4_o[7]~28 ));
defparam \u0_m0_wo0_mtree_add0_4_o[7]~27 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_4_o[7]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_4_o[8]~29 (
	.dataa(\u0_m0_wo0_mtree_mult1_8_sub_1_o[8]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_9_add_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_4_o[7]~28 ),
	.combout(\u0_m0_wo0_mtree_add0_4_o[8]~29_combout ),
	.cout(\u0_m0_wo0_mtree_add0_4_o[8]~30 ));
defparam \u0_m0_wo0_mtree_add0_4_o[8]~29 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_4_o[8]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_4_o[9]~31 (
	.dataa(\u0_m0_wo0_mtree_mult1_8_sub_1_o[9]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_9_add_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_4_o[8]~30 ),
	.combout(\u0_m0_wo0_mtree_add0_4_o[9]~31_combout ),
	.cout(\u0_m0_wo0_mtree_add0_4_o[9]~32 ));
defparam \u0_m0_wo0_mtree_add0_4_o[9]~31 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_4_o[9]~31 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add0_4_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_4_o[9]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_4_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_4_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_4_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_0_o[1]~12 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][0]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[1]~12_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[1]~13 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[1]~12 .lut_mask = 16'h6611;
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[1]~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_0_o[2]~14 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_0_o[1]~13 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[2]~14_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[2]~15 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[2]~14 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[2]~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_0_o[3]~16 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_0_o[2]~15 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[3]~16_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[3]~17 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[3]~16 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[3]~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_0_o[4]~18 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_0_o[3]~17 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[4]~18_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[4]~19 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[4]~18 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[4]~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_0_o[5]~20 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_0_o[4]~19 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[5]~20_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[5]~21 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[5]~20 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[5]~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_0_o[6]~22 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_0_o[5]~21 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[6]~22_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[6]~23 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[6]~22 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[6]~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_0_o[7]~24 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_0_o[6]~23 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[7]~24_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[7]~25 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[7]~24 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[7]~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_0_o[8]~26 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_0_o[7]~25 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[8]~26_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[8]~27 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[8]~26 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[8]~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_0_o[9]~28 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_0_o[8]~27 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[9]~28_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[9]~29 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[9]~28 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[9]~28 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_0_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_0_o[9]~28_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_0_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_0_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_0_o[8]~26_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_0_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_0_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_0_o[7]~24_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_0_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_0_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_0_o[6]~22_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_0_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_0_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_0_o[5]~20_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_0_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_0_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_0_o[4]~18_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_0_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_0_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_0_o[3]~16_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_0_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_0_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_0_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_0_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_0_o[2]~14_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_0_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[2] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_2_o[2]~13 (
	.dataa(\u0_m0_wo0_mtree_mult1_10_sub_0_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_0_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[2]~13_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[2]~14 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[2]~13 .lut_mask = 16'h66DD;
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[2]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_2_o[3]~15 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][1]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_0_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_2_o[2]~14 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[3]~15_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[3]~16 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[3]~15 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[3]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_2_o[4]~17 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][2]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_0_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_2_o[3]~16 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[4]~17_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[4]~18 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[4]~17 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[4]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_2_o[5]~19 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][3]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_0_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_2_o[4]~18 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[5]~19_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[5]~20 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[5]~19 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[5]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_2_o[6]~21 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][4]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_0_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_2_o[5]~20 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[6]~21_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[6]~22 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[6]~21 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[6]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_2_o[7]~23 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][5]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_0_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_2_o[6]~22 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[7]~23_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[7]~24 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[7]~23 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[7]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_2_o[8]~25 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][6]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_0_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_2_o[7]~24 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[8]~25_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[8]~26 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[8]~25 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[8]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_2_o[9]~27 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][7]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_0_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_2_o[8]~26 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[9]~27_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[9]~28 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[9]~27 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[9]~27 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_2_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_2_o[9]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_2_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_4_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_4_o[8]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_4_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_4_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_4_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_2_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_2_o[8]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_2_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_4_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_4_o[7]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_4_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_4_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_4_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_2_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_2_o[7]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_2_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_4_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_4_o[6]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_4_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_4_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_4_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_2_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_2_o[6]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_2_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_4_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_4_o[5]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_4_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_4_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_4_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_2_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_2_o[5]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_2_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_4_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_4_o[4]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_4_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_4_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_4_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_2_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_2_o[4]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_2_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_4_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_4_o[3]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_4_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_4_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_4_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_2_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_2_o[3]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_2_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_4_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_4_o[2]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_4_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_4_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_4_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_2_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_2_o[2]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_2_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_4_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_4_o[1]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_4_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_4_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_4_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_0_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_0_o[1]~12_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_0_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_2_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_0_o[1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_2_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_8_sub_1_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_8_sub_1_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_4_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_8_sub_1_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_4_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_4_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_4_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_2_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_0_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_2_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_2_o[0]~17 (
	.dataa(\u0_m0_wo0_mtree_add0_4_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_2_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_add1_2_o[0]~17_combout ),
	.cout(\u0_m0_wo0_mtree_add1_2_o[0]~18 ));
defparam \u0_m0_wo0_mtree_add1_2_o[0]~17 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_add1_2_o[0]~17 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_2_o[1]~19 (
	.dataa(\u0_m0_wo0_mtree_add0_4_o[1]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_2_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_2_o[0]~18 ),
	.combout(\u0_m0_wo0_mtree_add1_2_o[1]~19_combout ),
	.cout(\u0_m0_wo0_mtree_add1_2_o[1]~20 ));
defparam \u0_m0_wo0_mtree_add1_2_o[1]~19 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_2_o[1]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_2_o[2]~21 (
	.dataa(\u0_m0_wo0_mtree_add0_4_o[2]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_2_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_2_o[1]~20 ),
	.combout(\u0_m0_wo0_mtree_add1_2_o[2]~21_combout ),
	.cout(\u0_m0_wo0_mtree_add1_2_o[2]~22 ));
defparam \u0_m0_wo0_mtree_add1_2_o[2]~21 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_2_o[2]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_2_o[3]~23 (
	.dataa(\u0_m0_wo0_mtree_add0_4_o[3]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_2_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_2_o[2]~22 ),
	.combout(\u0_m0_wo0_mtree_add1_2_o[3]~23_combout ),
	.cout(\u0_m0_wo0_mtree_add1_2_o[3]~24 ));
defparam \u0_m0_wo0_mtree_add1_2_o[3]~23 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_2_o[3]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_2_o[4]~25 (
	.dataa(\u0_m0_wo0_mtree_add0_4_o[4]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_2_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_2_o[3]~24 ),
	.combout(\u0_m0_wo0_mtree_add1_2_o[4]~25_combout ),
	.cout(\u0_m0_wo0_mtree_add1_2_o[4]~26 ));
defparam \u0_m0_wo0_mtree_add1_2_o[4]~25 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_2_o[4]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_2_o[5]~27 (
	.dataa(\u0_m0_wo0_mtree_add0_4_o[5]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_2_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_2_o[4]~26 ),
	.combout(\u0_m0_wo0_mtree_add1_2_o[5]~27_combout ),
	.cout(\u0_m0_wo0_mtree_add1_2_o[5]~28 ));
defparam \u0_m0_wo0_mtree_add1_2_o[5]~27 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_2_o[5]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_2_o[6]~29 (
	.dataa(\u0_m0_wo0_mtree_add0_4_o[6]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_2_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_2_o[5]~28 ),
	.combout(\u0_m0_wo0_mtree_add1_2_o[6]~29_combout ),
	.cout(\u0_m0_wo0_mtree_add1_2_o[6]~30 ));
defparam \u0_m0_wo0_mtree_add1_2_o[6]~29 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_2_o[6]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_2_o[7]~31 (
	.dataa(\u0_m0_wo0_mtree_add0_4_o[7]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_2_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_2_o[6]~30 ),
	.combout(\u0_m0_wo0_mtree_add1_2_o[7]~31_combout ),
	.cout(\u0_m0_wo0_mtree_add1_2_o[7]~32 ));
defparam \u0_m0_wo0_mtree_add1_2_o[7]~31 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_2_o[7]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_2_o[8]~33 (
	.dataa(\u0_m0_wo0_mtree_add0_4_o[8]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_2_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_2_o[7]~32 ),
	.combout(\u0_m0_wo0_mtree_add1_2_o[8]~33_combout ),
	.cout(\u0_m0_wo0_mtree_add1_2_o[8]~34 ));
defparam \u0_m0_wo0_mtree_add1_2_o[8]~33 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_2_o[8]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_2_o[9]~35 (
	.dataa(\u0_m0_wo0_mtree_add0_4_o[9]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_2_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_2_o[8]~34 ),
	.combout(\u0_m0_wo0_mtree_add1_2_o[9]~35_combout ),
	.cout(\u0_m0_wo0_mtree_add1_2_o[9]~36 ));
defparam \u0_m0_wo0_mtree_add1_2_o[9]~35 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_2_o[9]~35 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add1_2_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_2_o[9]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_2_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_2_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_2_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_1_o[1]~13 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][0]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_1_o[1]~13_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_1_o[1]~14 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[1]~13 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[1]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_1_o[2]~15 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][2]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_1_o[1]~14 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_1_o[2]~15_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_1_o[2]~16 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[2]~15 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[2]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_1_o[3]~17 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][2]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_1_o[2]~16 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_1_o[3]~17_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_1_o[3]~18 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[3]~17 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[3]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_1_o[4]~19 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][4]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_1_o[3]~18 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_1_o[4]~19_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_1_o[4]~20 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[4]~19 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[4]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_1_o[5]~21 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][4]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_1_o[4]~20 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_1_o[5]~21_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_1_o[5]~22 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[5]~21 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[5]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_1_o[6]~23 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][6]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_1_o[5]~22 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_1_o[6]~23_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_1_o[6]~24 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[6]~23 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[6]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_1_o[7]~25 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][6]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_1_o[6]~24 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_1_o[7]~25_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_1_o[7]~26 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[7]~25 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[7]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_1_o[8]~27 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][8]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_1_o[7]~26 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_1_o[8]~27_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_1_o[8]~28 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[8]~27 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[8]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_1_o[9]~29 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][8]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_1_o[8]~28 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_1_o[9]~29_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_1_o[9]~30 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[9]~29 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[9]~29 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_12_add_1_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_1_o[9]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_1_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_1_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_1_o[8]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_1_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_1_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_1_o[7]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_1_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_1_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_1_o[6]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_1_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_1_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_1_o[5]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_1_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_1_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_1_o[4]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_1_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_1_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_1_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_1_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_1_o[3]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_1_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[3] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_3_o[3]~13 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_1_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_12_add_1_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_3_o[3]~13_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_3_o[3]~14 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[3]~13 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[3]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_3_o[4]~15 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][1]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_12_add_1_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_3_o[3]~14 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_3_o[4]~15_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_3_o[4]~16 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[4]~15 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[4]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_3_o[5]~17 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][2]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_12_add_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_3_o[4]~16 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_3_o[5]~17_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_3_o[5]~18 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[5]~17 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[5]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_3_o[6]~19 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][3]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_12_add_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_3_o[5]~18 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_3_o[6]~19_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_3_o[6]~20 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[6]~19 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[6]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_3_o[7]~21 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][4]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_12_add_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_3_o[6]~20 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_3_o[7]~21_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_3_o[7]~22 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[7]~21 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[7]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_3_o[8]~23 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][5]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_12_add_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_3_o[7]~22 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_3_o[8]~23_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_3_o[8]~24 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[8]~23 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[8]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_3_o[9]~25 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][6]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_12_add_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_3_o[8]~24 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_3_o[9]~25_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_3_o[9]~26 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[9]~25 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[9]~25 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_12_add_3_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_3_o[9]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_3_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_1_o[1]~15 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][0]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[1]~15_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[1]~16 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[1]~15 .lut_mask = 16'h6611;
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[1]~15 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_1_o[2]~17 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_1_o[1]~16 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[2]~17_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[2]~18 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[2]~17 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[2]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_1_o[3]~19 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][0]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_1_o[2]~18 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[3]~19_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[3]~20 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[3]~19 .lut_mask = 16'h962B;
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[3]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_1_o[4]~21 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][1]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_1_o[3]~20 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[4]~21_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[4]~22 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[4]~21 .lut_mask = 16'h694D;
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[4]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_1_o[5]~23 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][2]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_1_o[4]~22 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[5]~23_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[5]~24 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[5]~23 .lut_mask = 16'h962B;
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[5]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_1_o[6]~25 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][3]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_1_o[5]~24 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[6]~25_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[6]~26 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[6]~25 .lut_mask = 16'h694D;
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[6]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_1_o[7]~27 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][4]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_1_o[6]~26 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[7]~27_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[7]~28 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[7]~27 .lut_mask = 16'h962B;
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[7]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_1_o[8]~29 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][5]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_1_o[7]~28 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[8]~29_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[8]~30 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[8]~29 .lut_mask = 16'h694D;
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[8]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_1_o[9]~31 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][6]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_1_o[8]~30 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[9]~31_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[9]~32 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[9]~31 .lut_mask = 16'h962B;
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[9]~31 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_1_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[9]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_1_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_1_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[8]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_1_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_1_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[7]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_1_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_1_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[6]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_1_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_1_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_1_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_1_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[5]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_1_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[5] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_3_o[5]~13 (
	.dataa(\u0_m0_wo0_mtree_mult1_13_sub_1_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[5]~13_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[5]~14 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[5]~13 .lut_mask = 16'h66DD;
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[5]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_3_o[6]~15 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][1]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_3_o[5]~14 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[6]~15_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[6]~16 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[6]~15 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[6]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_3_o[7]~17 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][2]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_3_o[6]~16 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[7]~17_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[7]~18 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[7]~17 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[7]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_3_o[8]~19 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][3]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_3_o[7]~18 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[8]~19_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[8]~20 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[8]~19 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[8]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_3_o[9]~21 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][4]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_3_o[8]~20 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[9]~21_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[9]~22 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[9]~21 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[9]~21 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_3_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_3_o[9]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_3_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_3_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_3_o[8]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_3_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_3_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_3_o[8]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_3_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_3_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_3_o[7]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_3_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_3_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_3_o[7]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_3_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_3_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_3_o[6]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_3_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_3_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_3_o[6]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_3_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_3_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_3_o[5]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_3_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_3_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_3_o[5]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_3_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_3_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_3_o[4]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_3_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_1_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[4]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_1_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_3_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[4]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_3_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_3_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_3_o[3]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_3_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_1_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[3]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_1_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_3_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[3]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_3_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_1_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_1_o[2]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_1_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_3_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_1_o[2]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_3_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_1_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[2]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_1_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_3_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[2]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_3_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_1_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_1_o[1]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_1_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_3_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_1_o[1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_3_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_1_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[1]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_1_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_3_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_3_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_3_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_1_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_3_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_3_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_3_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_6_o[0]~19 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_3_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_3_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_add0_6_o[0]~19_combout ),
	.cout(\u0_m0_wo0_mtree_add0_6_o[0]~20 ));
defparam \u0_m0_wo0_mtree_add0_6_o[0]~19 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_add0_6_o[0]~19 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_6_o[1]~21 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_3_o[1]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_3_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_6_o[0]~20 ),
	.combout(\u0_m0_wo0_mtree_add0_6_o[1]~21_combout ),
	.cout(\u0_m0_wo0_mtree_add0_6_o[1]~22 ));
defparam \u0_m0_wo0_mtree_add0_6_o[1]~21 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_6_o[1]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_6_o[2]~23 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_3_o[2]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_3_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_6_o[1]~22 ),
	.combout(\u0_m0_wo0_mtree_add0_6_o[2]~23_combout ),
	.cout(\u0_m0_wo0_mtree_add0_6_o[2]~24 ));
defparam \u0_m0_wo0_mtree_add0_6_o[2]~23 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_6_o[2]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_6_o[3]~25 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_3_o[3]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_3_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_6_o[2]~24 ),
	.combout(\u0_m0_wo0_mtree_add0_6_o[3]~25_combout ),
	.cout(\u0_m0_wo0_mtree_add0_6_o[3]~26 ));
defparam \u0_m0_wo0_mtree_add0_6_o[3]~25 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_6_o[3]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_6_o[4]~27 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_3_o[4]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_3_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_6_o[3]~26 ),
	.combout(\u0_m0_wo0_mtree_add0_6_o[4]~27_combout ),
	.cout(\u0_m0_wo0_mtree_add0_6_o[4]~28 ));
defparam \u0_m0_wo0_mtree_add0_6_o[4]~27 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_6_o[4]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_6_o[5]~29 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_3_o[5]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_3_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_6_o[4]~28 ),
	.combout(\u0_m0_wo0_mtree_add0_6_o[5]~29_combout ),
	.cout(\u0_m0_wo0_mtree_add0_6_o[5]~30 ));
defparam \u0_m0_wo0_mtree_add0_6_o[5]~29 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_6_o[5]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_6_o[6]~31 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_3_o[6]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_3_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_6_o[5]~30 ),
	.combout(\u0_m0_wo0_mtree_add0_6_o[6]~31_combout ),
	.cout(\u0_m0_wo0_mtree_add0_6_o[6]~32 ));
defparam \u0_m0_wo0_mtree_add0_6_o[6]~31 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_6_o[6]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_6_o[7]~33 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_3_o[7]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_3_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_6_o[6]~32 ),
	.combout(\u0_m0_wo0_mtree_add0_6_o[7]~33_combout ),
	.cout(\u0_m0_wo0_mtree_add0_6_o[7]~34 ));
defparam \u0_m0_wo0_mtree_add0_6_o[7]~33 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_6_o[7]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_6_o[8]~35 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_3_o[8]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_3_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_6_o[7]~34 ),
	.combout(\u0_m0_wo0_mtree_add0_6_o[8]~35_combout ),
	.cout(\u0_m0_wo0_mtree_add0_6_o[8]~36 ));
defparam \u0_m0_wo0_mtree_add0_6_o[8]~35 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_6_o[8]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_6_o[9]~37 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_3_o[9]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_3_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_6_o[8]~36 ),
	.combout(\u0_m0_wo0_mtree_add0_6_o[9]~37_combout ),
	.cout(\u0_m0_wo0_mtree_add0_6_o[9]~38 ));
defparam \u0_m0_wo0_mtree_add0_6_o[9]~37 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_6_o[9]~37 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add0_6_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_6_o[9]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_6_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_6_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_6_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_1_o[2]~13 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][0]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_1_o[2]~13_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_1_o[2]~14 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[2]~13 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[2]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_1_o[3]~15 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][1]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_1_o[2]~14 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_1_o[3]~15_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_1_o[3]~16 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[3]~15 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[3]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_1_o[4]~17 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][2]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_1_o[3]~16 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_1_o[4]~17_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_1_o[4]~18 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[4]~17 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[4]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_1_o[5]~19 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][3]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_1_o[4]~18 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_1_o[5]~19_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_1_o[5]~20 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[5]~19 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[5]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_1_o[6]~21 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][4]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_1_o[5]~20 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_1_o[6]~21_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_1_o[6]~22 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[6]~21 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[6]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_1_o[7]~23 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][5]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_1_o[6]~22 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_1_o[7]~23_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_1_o[7]~24 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[7]~23 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[7]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_1_o[8]~25 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][6]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_1_o[7]~24 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_1_o[8]~25_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_1_o[8]~26 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[8]~25 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[8]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_1_o[9]~27 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][7]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_1_o[8]~26 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_1_o[9]~27_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_1_o[9]~28 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[9]~27 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[9]~27 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_14_add_1_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_1_o[9]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_1_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_1_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_1_o[8]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_1_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_1_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_1_o[7]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_1_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_1_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_1_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_1_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_1_o[6]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_1_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_1_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_1_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_1_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_1_o[5]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_1_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[5] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_3_o[5]~13 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_1_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_14_add_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_3_o[5]~13_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_3_o[5]~14 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[5]~13 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[5]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_3_o[6]~15 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_1_o[1]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_14_add_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_3_o[5]~14 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_3_o[6]~15_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_3_o[6]~16 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[6]~15 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[6]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_3_o[7]~17 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][2]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_14_add_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_3_o[6]~16 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_3_o[7]~17_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_3_o[7]~18 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[7]~17 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[7]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_3_o[8]~19 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][3]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_14_add_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_3_o[7]~18 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_3_o[8]~19_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_3_o[8]~20 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[8]~19 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[8]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_3_o[9]~21 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][4]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_14_add_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_3_o[8]~20 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_3_o[9]~21_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_3_o[9]~22 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[9]~21 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[9]~21 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_14_add_3_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_3_o[9]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_3_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_15_sub_1_o[1]~19 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][0]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[1]~19_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[1]~20 ));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[1]~19 .lut_mask = 16'h6611;
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[1]~19 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_15_sub_1_o[2]~21 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_15_sub_1_o[1]~20 ),
	.combout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[2]~21_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[2]~22 ));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[2]~21 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[2]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_15_sub_1_o[3]~23 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_15_sub_1_o[2]~22 ),
	.combout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[3]~23_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[3]~24 ));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[3]~23 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[3]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_15_sub_1_o[4]~25 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_15_sub_1_o[3]~24 ),
	.combout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[4]~25_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[4]~26 ));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[4]~25 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[4]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_15_sub_1_o[5]~27 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_15_sub_1_o[4]~26 ),
	.combout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[5]~27_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[5]~28 ));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[5]~27 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[5]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_15_sub_1_o[6]~29 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_15_sub_1_o[5]~28 ),
	.combout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[6]~29_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[6]~30 ));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[6]~29 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[6]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_15_sub_1_o[7]~31 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][0]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_15_sub_1_o[6]~30 ),
	.combout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[7]~31_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[7]~32 ));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[7]~31 .lut_mask = 16'h962B;
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[7]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_15_sub_1_o[8]~33 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][1]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_15_sub_1_o[7]~32 ),
	.combout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[8]~33_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[8]~34 ));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[8]~33 .lut_mask = 16'h694D;
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[8]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_15_sub_1_o[9]~35 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][2]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_15_sub_1_o[8]~34 ),
	.combout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[9]~35_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[9]~36 ));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[9]~35 .lut_mask = 16'h962B;
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[9]~35 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_15_sub_1_o[9]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_3_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_3_o[8]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_3_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_15_sub_1_o[8]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_3_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_3_o[7]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_3_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_15_sub_1_o[7]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_3_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_3_o[6]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_3_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_15_sub_1_o[6]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_3_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_3_o[5]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_3_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_15_sub_1_o[5]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_1_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_1_o[4]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_1_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_3_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_1_o[4]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_3_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_15_sub_1_o[4]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_1_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_1_o[3]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_1_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_3_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_1_o[3]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_3_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_15_sub_1_o[3]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_1_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_1_o[2]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_1_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_3_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_1_o[2]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_3_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_15_sub_1_o[2]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_3_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_1_o[1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_3_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_15_sub_1_o[1]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_3_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_1_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_3_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[0] (
	.clk(clk),
	.d(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[0]~21 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_add0_7_o[0]~21_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[0]~22 ));
defparam \u0_m0_wo0_mtree_add0_7_o[0]~21 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_add0_7_o[0]~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[1]~23 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[1]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_7_o[0]~22 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[1]~23_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[1]~24 ));
defparam \u0_m0_wo0_mtree_add0_7_o[1]~23 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_7_o[1]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[2]~25 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[2]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_7_o[1]~24 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[2]~25_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[2]~26 ));
defparam \u0_m0_wo0_mtree_add0_7_o[2]~25 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_7_o[2]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[3]~27 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[3]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_7_o[2]~26 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[3]~27_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[3]~28 ));
defparam \u0_m0_wo0_mtree_add0_7_o[3]~27 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_7_o[3]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[4]~29 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[4]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_7_o[3]~28 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[4]~29_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[4]~30 ));
defparam \u0_m0_wo0_mtree_add0_7_o[4]~29 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_7_o[4]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[5]~31 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[5]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_7_o[4]~30 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[5]~31_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[5]~32 ));
defparam \u0_m0_wo0_mtree_add0_7_o[5]~31 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_7_o[5]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[6]~33 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[6]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_7_o[5]~32 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[6]~33_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[6]~34 ));
defparam \u0_m0_wo0_mtree_add0_7_o[6]~33 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_7_o[6]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[7]~35 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[7]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_7_o[6]~34 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[7]~35_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[7]~36 ));
defparam \u0_m0_wo0_mtree_add0_7_o[7]~35 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_7_o[7]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[8]~37 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[8]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_7_o[7]~36 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[8]~37_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[8]~38 ));
defparam \u0_m0_wo0_mtree_add0_7_o[8]~37 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_7_o[8]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[9]~39 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[9]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_7_o[8]~38 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[9]~39_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[9]~40 ));
defparam \u0_m0_wo0_mtree_add0_7_o[9]~39 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_7_o[9]~39 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add0_7_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[9]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_6_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_6_o[8]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_6_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_6_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_6_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_7_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[8]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_6_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_6_o[7]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_6_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_6_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_6_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_7_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[7]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_6_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_6_o[6]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_6_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_6_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_6_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_7_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[6]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_6_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_6_o[5]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_6_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_6_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_6_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_7_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[5]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_6_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_6_o[4]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_6_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_6_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_6_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_7_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[4]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_6_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_6_o[3]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_6_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_6_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_6_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_7_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[3]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_6_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_6_o[2]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_6_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_6_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_6_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_7_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[2]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_6_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_6_o[1]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_6_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_6_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_6_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_7_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[1]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_6_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_6_o[0]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_6_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_6_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_6_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_7_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[0]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[0]~21 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_add1_3_o[0]~21_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[0]~22 ));
defparam \u0_m0_wo0_mtree_add1_3_o[0]~21 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_add1_3_o[0]~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[1]~23 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[1]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_3_o[0]~22 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[1]~23_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[1]~24 ));
defparam \u0_m0_wo0_mtree_add1_3_o[1]~23 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_3_o[1]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[2]~25 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[2]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_3_o[1]~24 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[2]~25_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[2]~26 ));
defparam \u0_m0_wo0_mtree_add1_3_o[2]~25 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_3_o[2]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[3]~27 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[3]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_3_o[2]~26 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[3]~27_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[3]~28 ));
defparam \u0_m0_wo0_mtree_add1_3_o[3]~27 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_3_o[3]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[4]~29 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[4]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_3_o[3]~28 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[4]~29_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[4]~30 ));
defparam \u0_m0_wo0_mtree_add1_3_o[4]~29 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_3_o[4]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[5]~31 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[5]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_3_o[4]~30 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[5]~31_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[5]~32 ));
defparam \u0_m0_wo0_mtree_add1_3_o[5]~31 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_3_o[5]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[6]~33 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[6]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_3_o[5]~32 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[6]~33_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[6]~34 ));
defparam \u0_m0_wo0_mtree_add1_3_o[6]~33 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_3_o[6]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[7]~35 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[7]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_3_o[6]~34 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[7]~35_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[7]~36 ));
defparam \u0_m0_wo0_mtree_add1_3_o[7]~35 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_3_o[7]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[8]~37 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[8]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_3_o[7]~36 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[8]~37_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[8]~38 ));
defparam \u0_m0_wo0_mtree_add1_3_o[8]~37 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_3_o[8]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[9]~39 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[9]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_3_o[8]~38 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[9]~39_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[9]~40 ));
defparam \u0_m0_wo0_mtree_add1_3_o[9]~39 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_3_o[9]~39 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add1_3_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[9]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_2_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_2_o[8]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_2_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_2_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_2_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_3_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[8]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_2_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_2_o[7]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_2_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_2_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_2_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_3_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[7]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_2_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_2_o[6]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_2_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_2_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_2_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_3_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[6]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_2_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_2_o[5]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_2_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_2_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_2_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_3_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[5]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_2_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_2_o[4]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_2_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_2_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_2_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_3_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[4]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_2_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_2_o[3]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_2_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_2_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_2_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_3_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[3]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_2_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_2_o[2]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_2_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_2_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_2_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_3_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[2]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_2_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_2_o[1]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_2_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_2_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_2_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_3_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[1]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_2_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_2_o[0]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_2_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_2_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_2_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_3_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[0]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[0]~21 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_add2_1_o[0]~21_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[0]~22 ));
defparam \u0_m0_wo0_mtree_add2_1_o[0]~21 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_add2_1_o[0]~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[1]~23 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[1]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_1_o[0]~22 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[1]~23_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[1]~24 ));
defparam \u0_m0_wo0_mtree_add2_1_o[1]~23 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_1_o[1]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[2]~25 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[2]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_1_o[1]~24 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[2]~25_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[2]~26 ));
defparam \u0_m0_wo0_mtree_add2_1_o[2]~25 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add2_1_o[2]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[3]~27 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[3]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_1_o[2]~26 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[3]~27_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[3]~28 ));
defparam \u0_m0_wo0_mtree_add2_1_o[3]~27 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_1_o[3]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[4]~29 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[4]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_1_o[3]~28 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[4]~29_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[4]~30 ));
defparam \u0_m0_wo0_mtree_add2_1_o[4]~29 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add2_1_o[4]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[5]~31 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[5]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_1_o[4]~30 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[5]~31_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[5]~32 ));
defparam \u0_m0_wo0_mtree_add2_1_o[5]~31 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_1_o[5]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[6]~33 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[6]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_1_o[5]~32 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[6]~33_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[6]~34 ));
defparam \u0_m0_wo0_mtree_add2_1_o[6]~33 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add2_1_o[6]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[7]~35 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[7]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_1_o[6]~34 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[7]~35_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[7]~36 ));
defparam \u0_m0_wo0_mtree_add2_1_o[7]~35 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_1_o[7]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[8]~37 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[8]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_1_o[7]~36 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[8]~37_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[8]~38 ));
defparam \u0_m0_wo0_mtree_add2_1_o[8]~37 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add2_1_o[8]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[9]~39 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[9]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_1_o[8]~38 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[9]~39_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[9]~40 ));
defparam \u0_m0_wo0_mtree_add2_1_o[9]~39 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_1_o[9]~39 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add2_1_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[9]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_1_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_1_o[8]~30_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_1_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_1_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_1_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_1_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[8]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_1_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_1_o[7]~28_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_1_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_1_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_1_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_1_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[7]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_1_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_1_o[6]~26_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_1_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_1_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_1_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_1_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[6]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_1_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_1_o[5]~24_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_1_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_1_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_1_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_1_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[5]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_1_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_1_o[4]~22_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_1_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_1_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_1_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_1_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[4]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_1_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_1_o[3]~20_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_1_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_1_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_1_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_1_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[3]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_1_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_1_o[2]~18_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_1_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_1_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_1_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_1_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[2]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_1_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_1_o[1]~16_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_1_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_1_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_1_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_1_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[1]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_1_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_1_o[0]~14_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_1_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_1_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_1_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_1_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[0]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[0]~21 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_add3_0_o[0]~21_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[0]~22 ));
defparam \u0_m0_wo0_mtree_add3_0_o[0]~21 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_add3_0_o[0]~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[1]~23 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[1]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_0_o[0]~22 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[1]~23_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[1]~24 ));
defparam \u0_m0_wo0_mtree_add3_0_o[1]~23 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_0_o[1]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[2]~25 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[2]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_0_o[1]~24 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[2]~25_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[2]~26 ));
defparam \u0_m0_wo0_mtree_add3_0_o[2]~25 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add3_0_o[2]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[3]~27 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[3]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_0_o[2]~26 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[3]~27_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[3]~28 ));
defparam \u0_m0_wo0_mtree_add3_0_o[3]~27 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_0_o[3]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[4]~29 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[4]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_0_o[3]~28 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[4]~29_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[4]~30 ));
defparam \u0_m0_wo0_mtree_add3_0_o[4]~29 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add3_0_o[4]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[5]~31 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[5]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_0_o[4]~30 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[5]~31_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[5]~32 ));
defparam \u0_m0_wo0_mtree_add3_0_o[5]~31 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_0_o[5]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[6]~33 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[6]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_0_o[5]~32 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[6]~33_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[6]~34 ));
defparam \u0_m0_wo0_mtree_add3_0_o[6]~33 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add3_0_o[6]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[7]~35 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[7]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_0_o[6]~34 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[7]~35_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[7]~36 ));
defparam \u0_m0_wo0_mtree_add3_0_o[7]~35 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_0_o[7]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[8]~37 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[8]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_0_o[7]~36 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[8]~37_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[8]~38 ));
defparam \u0_m0_wo0_mtree_add3_0_o[8]~37 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add3_0_o[8]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[9]~39 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[9]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_0_o[8]~38 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[9]~39_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[9]~40 ));
defparam \u0_m0_wo0_mtree_add3_0_o[9]~39 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_0_o[9]~39 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add3_0_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[9]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_1_o[2]~13 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][0]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_1_o[2]~13_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_1_o[2]~14 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[2]~13 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[2]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_1_o[3]~15 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][1]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_1_o[2]~14 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_1_o[3]~15_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_1_o[3]~16 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[3]~15 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[3]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_1_o[4]~17 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][2]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_1_o[3]~16 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_1_o[4]~17_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_1_o[4]~18 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[4]~17 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[4]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_1_o[5]~19 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][3]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_1_o[4]~18 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_1_o[5]~19_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_1_o[5]~20 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[5]~19 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[5]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_1_o[6]~21 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][4]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_1_o[5]~20 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_1_o[6]~21_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_1_o[6]~22 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[6]~21 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[6]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_1_o[7]~23 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][5]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_1_o[6]~22 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_1_o[7]~23_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_1_o[7]~24 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[7]~23 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[7]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_1_o[8]~25 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][6]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_1_o[7]~24 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_1_o[8]~25_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_1_o[8]~26 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[8]~25 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[8]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_1_o[9]~27 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][7]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_1_o[8]~26 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_1_o[9]~27_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_1_o[9]~28 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[9]~27 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[9]~27 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_16_add_1_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_1_o[9]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_1_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_1_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_1_o[8]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_1_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_1_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_1_o[7]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_1_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_1_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_1_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_1_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_1_o[6]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_1_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_1_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_1_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_1_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_1_o[5]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_1_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[5] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_3_o[5]~13 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_1_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_16_add_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_3_o[5]~13_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_3_o[5]~14 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[5]~13 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[5]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_3_o[6]~15 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_1_o[1]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_16_add_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_3_o[5]~14 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_3_o[6]~15_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_3_o[6]~16 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[6]~15 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[6]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_3_o[7]~17 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][2]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_16_add_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_3_o[6]~16 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_3_o[7]~17_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_3_o[7]~18 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[7]~17 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[7]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_3_o[8]~19 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][3]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_16_add_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_3_o[7]~18 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_3_o[8]~19_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_3_o[8]~20 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[8]~19 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[8]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_3_o[9]~21 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][4]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_16_add_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_3_o[8]~20 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_3_o[9]~21_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_3_o[9]~22 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[9]~21 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[9]~21 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_16_add_3_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_3_o[9]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_3_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_1_o[1]~15 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][0]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[1]~15_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[1]~16 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[1]~15 .lut_mask = 16'h6611;
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[1]~15 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_1_o[2]~17 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_1_o[1]~16 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[2]~17_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[2]~18 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[2]~17 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[2]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_1_o[3]~19 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][0]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_1_o[2]~18 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[3]~19_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[3]~20 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[3]~19 .lut_mask = 16'h962B;
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[3]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_1_o[4]~21 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][1]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_1_o[3]~20 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[4]~21_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[4]~22 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[4]~21 .lut_mask = 16'h694D;
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[4]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_1_o[5]~23 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][2]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_1_o[4]~22 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[5]~23_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[5]~24 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[5]~23 .lut_mask = 16'h962B;
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[5]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_1_o[6]~25 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][3]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_1_o[5]~24 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[6]~25_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[6]~26 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[6]~25 .lut_mask = 16'h694D;
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[6]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_1_o[7]~27 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][4]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_1_o[6]~26 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[7]~27_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[7]~28 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[7]~27 .lut_mask = 16'h962B;
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[7]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_1_o[8]~29 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][5]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_1_o[7]~28 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[8]~29_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[8]~30 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[8]~29 .lut_mask = 16'h694D;
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[8]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_1_o[9]~31 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][6]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_1_o[8]~30 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[9]~31_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[9]~32 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[9]~31 .lut_mask = 16'h962B;
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[9]~31 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_1_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[9]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_1_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_1_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[8]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_1_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_1_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[7]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_1_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_1_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[6]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_1_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_1_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_1_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_1_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[5]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_1_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[5] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_3_o[5]~13 (
	.dataa(\u0_m0_wo0_mtree_mult1_17_sub_1_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[5]~13_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[5]~14 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[5]~13 .lut_mask = 16'h66DD;
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[5]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_3_o[6]~15 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][1]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_3_o[5]~14 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[6]~15_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[6]~16 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[6]~15 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[6]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_3_o[7]~17 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][2]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_3_o[6]~16 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[7]~17_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[7]~18 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[7]~17 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[7]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_3_o[8]~19 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][3]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_3_o[7]~18 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[8]~19_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[8]~20 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[8]~19 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[8]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_3_o[9]~21 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][4]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_3_o[8]~20 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[9]~21_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[9]~22 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[9]~21 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[9]~21 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_3_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_3_o[9]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_3_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_3_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_3_o[8]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_3_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_3_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_3_o[8]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_3_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_3_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_3_o[7]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_3_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_3_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_3_o[7]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_3_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_3_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_3_o[6]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_3_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_3_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_3_o[6]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_3_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_3_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_3_o[5]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_3_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_3_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_3_o[5]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_3_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_1_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_1_o[4]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_1_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_3_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_1_o[4]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_3_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_1_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[4]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_1_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_3_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[4]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_3_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_1_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_1_o[3]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_1_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_3_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_1_o[3]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_3_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_1_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[3]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_1_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_3_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[3]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_3_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_1_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_1_o[2]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_1_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_3_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_1_o[2]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_3_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_1_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[2]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_1_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_3_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[2]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_3_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_3_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_1_o[1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_3_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_1_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[1]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_1_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_3_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_3_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_3_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_1_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_3_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_3_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_3_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_8_o[0]~19 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_3_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_3_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_add0_8_o[0]~19_combout ),
	.cout(\u0_m0_wo0_mtree_add0_8_o[0]~20 ));
defparam \u0_m0_wo0_mtree_add0_8_o[0]~19 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_add0_8_o[0]~19 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_8_o[1]~21 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_3_o[1]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_3_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_8_o[0]~20 ),
	.combout(\u0_m0_wo0_mtree_add0_8_o[1]~21_combout ),
	.cout(\u0_m0_wo0_mtree_add0_8_o[1]~22 ));
defparam \u0_m0_wo0_mtree_add0_8_o[1]~21 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_8_o[1]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_8_o[2]~23 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_3_o[2]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_3_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_8_o[1]~22 ),
	.combout(\u0_m0_wo0_mtree_add0_8_o[2]~23_combout ),
	.cout(\u0_m0_wo0_mtree_add0_8_o[2]~24 ));
defparam \u0_m0_wo0_mtree_add0_8_o[2]~23 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_8_o[2]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_8_o[3]~25 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_3_o[3]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_3_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_8_o[2]~24 ),
	.combout(\u0_m0_wo0_mtree_add0_8_o[3]~25_combout ),
	.cout(\u0_m0_wo0_mtree_add0_8_o[3]~26 ));
defparam \u0_m0_wo0_mtree_add0_8_o[3]~25 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_8_o[3]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_8_o[4]~27 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_3_o[4]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_3_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_8_o[3]~26 ),
	.combout(\u0_m0_wo0_mtree_add0_8_o[4]~27_combout ),
	.cout(\u0_m0_wo0_mtree_add0_8_o[4]~28 ));
defparam \u0_m0_wo0_mtree_add0_8_o[4]~27 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_8_o[4]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_8_o[5]~29 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_3_o[5]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_3_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_8_o[4]~28 ),
	.combout(\u0_m0_wo0_mtree_add0_8_o[5]~29_combout ),
	.cout(\u0_m0_wo0_mtree_add0_8_o[5]~30 ));
defparam \u0_m0_wo0_mtree_add0_8_o[5]~29 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_8_o[5]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_8_o[6]~31 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_3_o[6]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_3_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_8_o[5]~30 ),
	.combout(\u0_m0_wo0_mtree_add0_8_o[6]~31_combout ),
	.cout(\u0_m0_wo0_mtree_add0_8_o[6]~32 ));
defparam \u0_m0_wo0_mtree_add0_8_o[6]~31 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_8_o[6]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_8_o[7]~33 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_3_o[7]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_3_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_8_o[6]~32 ),
	.combout(\u0_m0_wo0_mtree_add0_8_o[7]~33_combout ),
	.cout(\u0_m0_wo0_mtree_add0_8_o[7]~34 ));
defparam \u0_m0_wo0_mtree_add0_8_o[7]~33 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_8_o[7]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_8_o[8]~35 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_3_o[8]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_3_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_8_o[7]~34 ),
	.combout(\u0_m0_wo0_mtree_add0_8_o[8]~35_combout ),
	.cout(\u0_m0_wo0_mtree_add0_8_o[8]~36 ));
defparam \u0_m0_wo0_mtree_add0_8_o[8]~35 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_8_o[8]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_8_o[9]~37 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_3_o[9]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_3_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_8_o[8]~36 ),
	.combout(\u0_m0_wo0_mtree_add0_8_o[9]~37_combout ),
	.cout(\u0_m0_wo0_mtree_add0_8_o[9]~38 ));
defparam \u0_m0_wo0_mtree_add0_8_o[9]~37 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_8_o[9]~37 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add0_8_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_8_o[9]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_8_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_8_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_8_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_1_o[1]~13 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][0]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_1_o[1]~13_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_1_o[1]~14 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[1]~13 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[1]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_1_o[2]~15 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][2]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_1_o[1]~14 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_1_o[2]~15_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_1_o[2]~16 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[2]~15 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[2]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_1_o[3]~17 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][2]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_1_o[2]~16 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_1_o[3]~17_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_1_o[3]~18 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[3]~17 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[3]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_1_o[4]~19 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][4]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_1_o[3]~18 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_1_o[4]~19_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_1_o[4]~20 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[4]~19 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[4]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_1_o[5]~21 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][4]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_1_o[4]~20 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_1_o[5]~21_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_1_o[5]~22 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[5]~21 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[5]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_1_o[6]~23 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][6]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_1_o[5]~22 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_1_o[6]~23_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_1_o[6]~24 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[6]~23 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[6]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_1_o[7]~25 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][6]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_1_o[6]~24 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_1_o[7]~25_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_1_o[7]~26 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[7]~25 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[7]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_1_o[8]~27 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][8]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_1_o[7]~26 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_1_o[8]~27_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_1_o[8]~28 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[8]~27 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[8]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_1_o[9]~29 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][8]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_1_o[8]~28 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_1_o[9]~29_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_1_o[9]~30 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[9]~29 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[9]~29 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_18_add_1_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_1_o[9]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_1_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_1_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_1_o[8]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_1_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_1_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_1_o[7]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_1_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_1_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_1_o[6]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_1_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_1_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_1_o[5]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_1_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_1_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_1_o[4]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_1_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_1_o[0] (
	.clk(clk),
	.d(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_1_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_1_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_1_o[3]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_1_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[3] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_3_o[3]~13 (
	.dataa(\u0_m0_wo0_mtree_mult1_18_add_1_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_1_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_3_o[3]~13_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_3_o[3]~14 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[3]~13 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[3]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_3_o[4]~15 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][1]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_1_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_3_o[3]~14 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_3_o[4]~15_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_3_o[4]~16 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[4]~15 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[4]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_3_o[5]~17 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][2]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_3_o[4]~16 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_3_o[5]~17_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_3_o[5]~18 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[5]~17 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[5]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_3_o[6]~19 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][3]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_3_o[5]~18 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_3_o[6]~19_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_3_o[6]~20 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[6]~19 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[6]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_3_o[7]~21 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][4]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_3_o[6]~20 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_3_o[7]~21_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_3_o[7]~22 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[7]~21 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[7]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_3_o[8]~23 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][5]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_3_o[7]~22 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_3_o[8]~23_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_3_o[8]~24 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[8]~23 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[8]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_3_o[9]~25 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][6]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_3_o[8]~24 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_3_o[9]~25_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_3_o[9]~26 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[9]~25 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[9]~25 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_18_add_3_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_3_o[9]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_3_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_8_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_8_o[8]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_8_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_8_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_8_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_3_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_3_o[8]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_3_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_8_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_8_o[7]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_8_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_8_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_8_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_3_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_3_o[7]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_3_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_8_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_8_o[6]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_8_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_8_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_8_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_3_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_3_o[6]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_3_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_8_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_8_o[5]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_8_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_8_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_8_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_3_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_3_o[5]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_3_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_8_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_8_o[4]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_8_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_8_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_8_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_3_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_3_o[4]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_3_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_8_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_8_o[3]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_8_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_8_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_8_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_3_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_3_o[3]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_3_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_8_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_8_o[2]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_8_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_8_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_8_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_1_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_1_o[2]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_1_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_3_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_1_o[2]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_3_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_8_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_8_o[1]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_8_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_8_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_8_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_1_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_1_o[1]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_1_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_3_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_1_o[1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_3_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_8_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_8_o[0]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_8_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_8_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_8_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_3_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_1_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_3_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[0]~20 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_add1_4_o[0]~20_combout ),
	.cout(\u0_m0_wo0_mtree_add1_4_o[0]~21 ));
defparam \u0_m0_wo0_mtree_add1_4_o[0]~20 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_add1_4_o[0]~20 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[1]~22 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[1]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_4_o[0]~21 ),
	.combout(\u0_m0_wo0_mtree_add1_4_o[1]~22_combout ),
	.cout(\u0_m0_wo0_mtree_add1_4_o[1]~23 ));
defparam \u0_m0_wo0_mtree_add1_4_o[1]~22 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_4_o[1]~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[2]~24 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[2]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_4_o[1]~23 ),
	.combout(\u0_m0_wo0_mtree_add1_4_o[2]~24_combout ),
	.cout(\u0_m0_wo0_mtree_add1_4_o[2]~25 ));
defparam \u0_m0_wo0_mtree_add1_4_o[2]~24 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_4_o[2]~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[3]~26 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[3]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_4_o[2]~25 ),
	.combout(\u0_m0_wo0_mtree_add1_4_o[3]~26_combout ),
	.cout(\u0_m0_wo0_mtree_add1_4_o[3]~27 ));
defparam \u0_m0_wo0_mtree_add1_4_o[3]~26 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_4_o[3]~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[4]~28 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[4]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_4_o[3]~27 ),
	.combout(\u0_m0_wo0_mtree_add1_4_o[4]~28_combout ),
	.cout(\u0_m0_wo0_mtree_add1_4_o[4]~29 ));
defparam \u0_m0_wo0_mtree_add1_4_o[4]~28 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_4_o[4]~28 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[5]~30 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[5]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_4_o[4]~29 ),
	.combout(\u0_m0_wo0_mtree_add1_4_o[5]~30_combout ),
	.cout(\u0_m0_wo0_mtree_add1_4_o[5]~31 ));
defparam \u0_m0_wo0_mtree_add1_4_o[5]~30 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_4_o[5]~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[6]~32 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[6]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_4_o[5]~31 ),
	.combout(\u0_m0_wo0_mtree_add1_4_o[6]~32_combout ),
	.cout(\u0_m0_wo0_mtree_add1_4_o[6]~33 ));
defparam \u0_m0_wo0_mtree_add1_4_o[6]~32 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_4_o[6]~32 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[7]~34 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[7]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_4_o[6]~33 ),
	.combout(\u0_m0_wo0_mtree_add1_4_o[7]~34_combout ),
	.cout(\u0_m0_wo0_mtree_add1_4_o[7]~35 ));
defparam \u0_m0_wo0_mtree_add1_4_o[7]~34 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_4_o[7]~34 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[8]~36 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[8]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_4_o[7]~35 ),
	.combout(\u0_m0_wo0_mtree_add1_4_o[8]~36_combout ),
	.cout(\u0_m0_wo0_mtree_add1_4_o[8]~37 ));
defparam \u0_m0_wo0_mtree_add1_4_o[8]~36 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_4_o[8]~36 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[9]~38 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[9]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_4_o[8]~37 ),
	.combout(\u0_m0_wo0_mtree_add1_4_o[9]~38_combout ),
	.cout(\u0_m0_wo0_mtree_add1_4_o[9]~39 ));
defparam \u0_m0_wo0_mtree_add1_4_o[9]~38 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_4_o[9]~38 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add1_4_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[9]~38_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_0_o[1]~12 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][0]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[1]~12_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[1]~13 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[1]~12 .lut_mask = 16'h6611;
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[1]~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_0_o[2]~14 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_0_o[1]~13 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[2]~14_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[2]~15 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[2]~14 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[2]~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_0_o[3]~16 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_0_o[2]~15 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[3]~16_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[3]~17 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[3]~16 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[3]~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_0_o[4]~18 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_0_o[3]~17 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[4]~18_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[4]~19 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[4]~18 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[4]~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_0_o[5]~20 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_0_o[4]~19 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[5]~20_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[5]~21 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[5]~20 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[5]~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_0_o[6]~22 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_0_o[5]~21 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[6]~22_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[6]~23 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[6]~22 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[6]~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_0_o[7]~24 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_0_o[6]~23 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[7]~24_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[7]~25 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[7]~24 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[7]~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_0_o[8]~26 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_0_o[7]~25 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[8]~26_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[8]~27 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[8]~26 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[8]~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_0_o[9]~28 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_0_o[8]~27 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[9]~28_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[9]~29 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[9]~28 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[9]~28 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_0_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_0_o[9]~28_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_0_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_0_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_0_o[8]~26_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_0_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_0_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_0_o[7]~24_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_0_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_0_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_0_o[6]~22_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_0_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_0_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_0_o[5]~20_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_0_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_0_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_0_o[4]~18_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_0_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_0_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_0_o[3]~16_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_0_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_0_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_0_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_0_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_0_o[2]~14_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_0_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[2] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_2_o[2]~13 (
	.dataa(\u0_m0_wo0_mtree_mult1_20_sub_0_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_20_sub_0_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[2]~13_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[2]~14 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[2]~13 .lut_mask = 16'h66DD;
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[2]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_2_o[3]~15 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][1]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_20_sub_0_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_2_o[2]~14 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[3]~15_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[3]~16 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[3]~15 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[3]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_2_o[4]~17 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][2]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_20_sub_0_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_2_o[3]~16 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[4]~17_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[4]~18 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[4]~17 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[4]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_2_o[5]~19 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][3]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_20_sub_0_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_2_o[4]~18 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[5]~19_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[5]~20 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[5]~19 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[5]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_2_o[6]~21 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][4]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_20_sub_0_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_2_o[5]~20 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[6]~21_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[6]~22 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[6]~21 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[6]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_2_o[7]~23 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][5]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_20_sub_0_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_2_o[6]~22 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[7]~23_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[7]~24 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[7]~23 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[7]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_2_o[8]~25 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][6]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_20_sub_0_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_2_o[7]~24 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[8]~25_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[8]~26 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[8]~25 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[8]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_2_o[9]~27 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][7]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_20_sub_0_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_2_o[8]~26 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[9]~27_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[9]~28 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[9]~27 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[9]~27 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_2_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_2_o[9]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_2_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_21_add_1_o[1]~13 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][0]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_21_add_1_o[1]~13_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_21_add_1_o[1]~14 ));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[1]~13 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[1]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_21_add_1_o[2]~15 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][2]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_21_add_1_o[1]~14 ),
	.combout(\u0_m0_wo0_mtree_mult1_21_add_1_o[2]~15_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_21_add_1_o[2]~16 ));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[2]~15 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[2]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_21_add_1_o[3]~17 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][2]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_21_add_1_o[2]~16 ),
	.combout(\u0_m0_wo0_mtree_mult1_21_add_1_o[3]~17_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_21_add_1_o[3]~18 ));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[3]~17 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[3]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_21_add_1_o[4]~19 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][4]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_21_add_1_o[3]~18 ),
	.combout(\u0_m0_wo0_mtree_mult1_21_add_1_o[4]~19_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_21_add_1_o[4]~20 ));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[4]~19 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[4]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_21_add_1_o[5]~21 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][4]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_21_add_1_o[4]~20 ),
	.combout(\u0_m0_wo0_mtree_mult1_21_add_1_o[5]~21_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_21_add_1_o[5]~22 ));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[5]~21 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[5]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_21_add_1_o[6]~23 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][6]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_21_add_1_o[5]~22 ),
	.combout(\u0_m0_wo0_mtree_mult1_21_add_1_o[6]~23_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_21_add_1_o[6]~24 ));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[6]~23 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[6]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_21_add_1_o[7]~25 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][6]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_21_add_1_o[6]~24 ),
	.combout(\u0_m0_wo0_mtree_mult1_21_add_1_o[7]~25_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_21_add_1_o[7]~26 ));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[7]~25 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[7]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_21_add_1_o[8]~27 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][8]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_21_add_1_o[7]~26 ),
	.combout(\u0_m0_wo0_mtree_mult1_21_add_1_o[8]~27_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_21_add_1_o[8]~28 ));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[8]~27 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[8]~27 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_21_add_1_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_21_add_1_o[8]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_21_add_1_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_2_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_2_o[8]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_2_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_21_add_1_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_21_add_1_o[7]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_21_add_1_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_2_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_2_o[7]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_2_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_21_add_1_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_21_add_1_o[6]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_21_add_1_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_2_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_2_o[6]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_2_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_21_add_1_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_21_add_1_o[5]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_21_add_1_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_2_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_2_o[5]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_2_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_21_add_1_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_21_add_1_o[4]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_21_add_1_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_2_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_2_o[4]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_2_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_21_add_1_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_21_add_1_o[3]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_21_add_1_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_2_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_2_o[3]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_2_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_21_add_1_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_21_add_1_o[2]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_21_add_1_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_2_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_2_o[2]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_2_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_21_add_1_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_21_add_1_o[1]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_21_add_1_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_0_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_0_o[1]~12_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_0_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_2_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_0_o[1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_2_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_21_add_1_o[0] (
	.clk(clk),
	.d(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_21_add_1_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_10_o[1]~15 (
	.dataa(\u0_m0_wo0_mtree_mult1_20_sub_2_o[1]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_21_add_1_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_add0_10_o[1]~15_combout ),
	.cout(\u0_m0_wo0_mtree_add0_10_o[1]~16 ));
defparam \u0_m0_wo0_mtree_add0_10_o[1]~15 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_add0_10_o[1]~15 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_10_o[2]~17 (
	.dataa(\u0_m0_wo0_mtree_mult1_20_sub_2_o[2]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_21_add_1_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_10_o[1]~16 ),
	.combout(\u0_m0_wo0_mtree_add0_10_o[2]~17_combout ),
	.cout(\u0_m0_wo0_mtree_add0_10_o[2]~18 ));
defparam \u0_m0_wo0_mtree_add0_10_o[2]~17 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_10_o[2]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_10_o[3]~19 (
	.dataa(\u0_m0_wo0_mtree_mult1_20_sub_2_o[3]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_21_add_1_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_10_o[2]~18 ),
	.combout(\u0_m0_wo0_mtree_add0_10_o[3]~19_combout ),
	.cout(\u0_m0_wo0_mtree_add0_10_o[3]~20 ));
defparam \u0_m0_wo0_mtree_add0_10_o[3]~19 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_10_o[3]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_10_o[4]~21 (
	.dataa(\u0_m0_wo0_mtree_mult1_20_sub_2_o[4]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_21_add_1_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_10_o[3]~20 ),
	.combout(\u0_m0_wo0_mtree_add0_10_o[4]~21_combout ),
	.cout(\u0_m0_wo0_mtree_add0_10_o[4]~22 ));
defparam \u0_m0_wo0_mtree_add0_10_o[4]~21 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_10_o[4]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_10_o[5]~23 (
	.dataa(\u0_m0_wo0_mtree_mult1_20_sub_2_o[5]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_21_add_1_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_10_o[4]~22 ),
	.combout(\u0_m0_wo0_mtree_add0_10_o[5]~23_combout ),
	.cout(\u0_m0_wo0_mtree_add0_10_o[5]~24 ));
defparam \u0_m0_wo0_mtree_add0_10_o[5]~23 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_10_o[5]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_10_o[6]~25 (
	.dataa(\u0_m0_wo0_mtree_mult1_20_sub_2_o[6]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_21_add_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_10_o[5]~24 ),
	.combout(\u0_m0_wo0_mtree_add0_10_o[6]~25_combout ),
	.cout(\u0_m0_wo0_mtree_add0_10_o[6]~26 ));
defparam \u0_m0_wo0_mtree_add0_10_o[6]~25 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_10_o[6]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_10_o[7]~27 (
	.dataa(\u0_m0_wo0_mtree_mult1_20_sub_2_o[7]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_21_add_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_10_o[6]~26 ),
	.combout(\u0_m0_wo0_mtree_add0_10_o[7]~27_combout ),
	.cout(\u0_m0_wo0_mtree_add0_10_o[7]~28 ));
defparam \u0_m0_wo0_mtree_add0_10_o[7]~27 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_10_o[7]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_10_o[8]~29 (
	.dataa(\u0_m0_wo0_mtree_mult1_20_sub_2_o[8]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_21_add_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_10_o[7]~28 ),
	.combout(\u0_m0_wo0_mtree_add0_10_o[8]~29_combout ),
	.cout(\u0_m0_wo0_mtree_add0_10_o[8]~30 ));
defparam \u0_m0_wo0_mtree_add0_10_o[8]~29 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_10_o[8]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_10_o[9]~31 (
	.dataa(\u0_m0_wo0_mtree_mult1_20_sub_2_o[9]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_21_add_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_10_o[8]~30 ),
	.combout(\u0_m0_wo0_mtree_add0_10_o[9]~31_combout ),
	.cout(\u0_m0_wo0_mtree_add0_10_o[9]~32 ));
defparam \u0_m0_wo0_mtree_add0_10_o[9]~31 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_10_o[9]~31 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add0_10_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_10_o[9]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_10_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_10_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_10_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_22_sub_1_o[2]~13 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][0]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[2]~13_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[2]~14 ));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[2]~13 .lut_mask = 16'h66DD;
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[2]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_22_sub_1_o[3]~15 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][1]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_22_sub_1_o[2]~14 ),
	.combout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[3]~15_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[3]~16 ));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[3]~15 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[3]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_22_sub_1_o[4]~17 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][2]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_22_sub_1_o[3]~16 ),
	.combout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[4]~17_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[4]~18 ));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[4]~17 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[4]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_22_sub_1_o[5]~19 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][3]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_22_sub_1_o[4]~18 ),
	.combout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[5]~19_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[5]~20 ));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[5]~19 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[5]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_22_sub_1_o[6]~21 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][4]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_22_sub_1_o[5]~20 ),
	.combout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[6]~21_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[6]~22 ));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[6]~21 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[6]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_22_sub_1_o[7]~23 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][5]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_22_sub_1_o[6]~22 ),
	.combout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[7]~23_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[7]~24 ));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[7]~23 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[7]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_22_sub_1_o[8]~25 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][6]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_22_sub_1_o[7]~24 ),
	.combout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[8]~25_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[8]~26 ));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[8]~25 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[8]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_22_sub_1_o[9]~27 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][7]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_22_sub_1_o[8]~26 ),
	.combout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[9]~27_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[9]~28 ));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[9]~27 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[9]~27 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_22_sub_1_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_22_sub_1_o[9]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_22_sub_1_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_10_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_10_o[8]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_10_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_10_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_10_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_22_sub_1_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_22_sub_1_o[8]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_22_sub_1_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_10_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_10_o[7]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_10_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_10_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_10_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_22_sub_1_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_22_sub_1_o[7]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_22_sub_1_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_10_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_10_o[6]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_10_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_10_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_10_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_22_sub_1_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_22_sub_1_o[6]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_22_sub_1_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_10_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_10_o[5]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_10_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_10_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_10_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_22_sub_1_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_22_sub_1_o[5]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_22_sub_1_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_10_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_10_o[4]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_10_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_10_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_10_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_22_sub_1_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_22_sub_1_o[4]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_22_sub_1_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_10_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_10_o[3]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_10_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_10_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_10_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_22_sub_1_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_22_sub_1_o[3]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_22_sub_1_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_10_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_10_o[2]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_10_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_10_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_10_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_22_sub_1_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_22_sub_1_o[2]~13_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_22_sub_1_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_10_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_10_o[1]~15_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_10_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_10_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_10_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_22_sub_1_o[1] (
	.clk(clk),
	.d(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][1]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_22_sub_1_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_2_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_0_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_2_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_10_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_2_o[0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_10_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_10_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_10_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_22_sub_1_o[0] (
	.clk(clk),
	.d(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_22_sub_1_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_5_o[0]~17 (
	.dataa(\u0_m0_wo0_mtree_add0_10_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_22_sub_1_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_add1_5_o[0]~17_combout ),
	.cout(\u0_m0_wo0_mtree_add1_5_o[0]~18 ));
defparam \u0_m0_wo0_mtree_add1_5_o[0]~17 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_add1_5_o[0]~17 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_5_o[1]~19 (
	.dataa(\u0_m0_wo0_mtree_add0_10_o[1]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_22_sub_1_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_5_o[0]~18 ),
	.combout(\u0_m0_wo0_mtree_add1_5_o[1]~19_combout ),
	.cout(\u0_m0_wo0_mtree_add1_5_o[1]~20 ));
defparam \u0_m0_wo0_mtree_add1_5_o[1]~19 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_5_o[1]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_5_o[2]~21 (
	.dataa(\u0_m0_wo0_mtree_add0_10_o[2]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_22_sub_1_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_5_o[1]~20 ),
	.combout(\u0_m0_wo0_mtree_add1_5_o[2]~21_combout ),
	.cout(\u0_m0_wo0_mtree_add1_5_o[2]~22 ));
defparam \u0_m0_wo0_mtree_add1_5_o[2]~21 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_5_o[2]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_5_o[3]~23 (
	.dataa(\u0_m0_wo0_mtree_add0_10_o[3]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_22_sub_1_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_5_o[2]~22 ),
	.combout(\u0_m0_wo0_mtree_add1_5_o[3]~23_combout ),
	.cout(\u0_m0_wo0_mtree_add1_5_o[3]~24 ));
defparam \u0_m0_wo0_mtree_add1_5_o[3]~23 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_5_o[3]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_5_o[4]~25 (
	.dataa(\u0_m0_wo0_mtree_add0_10_o[4]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_22_sub_1_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_5_o[3]~24 ),
	.combout(\u0_m0_wo0_mtree_add1_5_o[4]~25_combout ),
	.cout(\u0_m0_wo0_mtree_add1_5_o[4]~26 ));
defparam \u0_m0_wo0_mtree_add1_5_o[4]~25 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_5_o[4]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_5_o[5]~27 (
	.dataa(\u0_m0_wo0_mtree_add0_10_o[5]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_22_sub_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_5_o[4]~26 ),
	.combout(\u0_m0_wo0_mtree_add1_5_o[5]~27_combout ),
	.cout(\u0_m0_wo0_mtree_add1_5_o[5]~28 ));
defparam \u0_m0_wo0_mtree_add1_5_o[5]~27 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_5_o[5]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_5_o[6]~29 (
	.dataa(\u0_m0_wo0_mtree_add0_10_o[6]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_22_sub_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_5_o[5]~28 ),
	.combout(\u0_m0_wo0_mtree_add1_5_o[6]~29_combout ),
	.cout(\u0_m0_wo0_mtree_add1_5_o[6]~30 ));
defparam \u0_m0_wo0_mtree_add1_5_o[6]~29 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_5_o[6]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_5_o[7]~31 (
	.dataa(\u0_m0_wo0_mtree_add0_10_o[7]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_22_sub_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_5_o[6]~30 ),
	.combout(\u0_m0_wo0_mtree_add1_5_o[7]~31_combout ),
	.cout(\u0_m0_wo0_mtree_add1_5_o[7]~32 ));
defparam \u0_m0_wo0_mtree_add1_5_o[7]~31 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_5_o[7]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_5_o[8]~33 (
	.dataa(\u0_m0_wo0_mtree_add0_10_o[8]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_22_sub_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_5_o[7]~32 ),
	.combout(\u0_m0_wo0_mtree_add1_5_o[8]~33_combout ),
	.cout(\u0_m0_wo0_mtree_add1_5_o[8]~34 ));
defparam \u0_m0_wo0_mtree_add1_5_o[8]~33 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_5_o[8]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_5_o[9]~35 (
	.dataa(\u0_m0_wo0_mtree_add0_10_o[9]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_22_sub_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_5_o[8]~34 ),
	.combout(\u0_m0_wo0_mtree_add1_5_o[9]~35_combout ),
	.cout(\u0_m0_wo0_mtree_add1_5_o[9]~36 ));
defparam \u0_m0_wo0_mtree_add1_5_o[9]~35 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_5_o[9]~35 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add1_5_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_5_o[9]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_5_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_5_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_5_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_4_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[8]~36_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_5_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_5_o[8]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_5_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_5_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_5_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_4_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[7]~34_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_5_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_5_o[7]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_5_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_5_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_5_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_4_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[6]~32_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_5_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_5_o[6]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_5_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_5_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_5_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_4_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[5]~30_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_5_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_5_o[5]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_5_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_5_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_5_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_4_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[4]~28_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_5_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_5_o[4]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_5_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_5_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_5_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_4_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[3]~26_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_5_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_5_o[3]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_5_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_5_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_5_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_4_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[2]~24_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_5_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_5_o[2]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_5_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_5_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_5_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_4_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[1]~22_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_5_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_5_o[1]~19_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_5_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_5_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_5_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_4_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[0]~20_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_5_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_5_o[0]~17_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_5_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_5_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_5_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[0]~21 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_add2_2_o[0]~21_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[0]~22 ));
defparam \u0_m0_wo0_mtree_add2_2_o[0]~21 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_add2_2_o[0]~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[1]~23 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[1]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_2_o[0]~22 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[1]~23_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[1]~24 ));
defparam \u0_m0_wo0_mtree_add2_2_o[1]~23 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_2_o[1]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[2]~25 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[2]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_2_o[1]~24 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[2]~25_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[2]~26 ));
defparam \u0_m0_wo0_mtree_add2_2_o[2]~25 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add2_2_o[2]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[3]~27 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[3]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_2_o[2]~26 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[3]~27_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[3]~28 ));
defparam \u0_m0_wo0_mtree_add2_2_o[3]~27 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_2_o[3]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[4]~29 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[4]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_2_o[3]~28 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[4]~29_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[4]~30 ));
defparam \u0_m0_wo0_mtree_add2_2_o[4]~29 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add2_2_o[4]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[5]~31 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[5]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_2_o[4]~30 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[5]~31_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[5]~32 ));
defparam \u0_m0_wo0_mtree_add2_2_o[5]~31 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_2_o[5]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[6]~33 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[6]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_2_o[5]~32 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[6]~33_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[6]~34 ));
defparam \u0_m0_wo0_mtree_add2_2_o[6]~33 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add2_2_o[6]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[7]~35 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[7]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_2_o[6]~34 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[7]~35_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[7]~36 ));
defparam \u0_m0_wo0_mtree_add2_2_o[7]~35 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_2_o[7]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[8]~37 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[8]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_2_o[7]~36 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[8]~37_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[8]~38 ));
defparam \u0_m0_wo0_mtree_add2_2_o[8]~37 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add2_2_o[8]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[9]~39 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[9]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_2_o[8]~38 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[9]~39_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[9]~40 ));
defparam \u0_m0_wo0_mtree_add2_2_o[9]~39 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_2_o[9]~39 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add2_2_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[9]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_25_sub_0_o[1]~12 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][0]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[1]~12_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[1]~13 ));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[1]~12 .lut_mask = 16'h6611;
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[1]~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_25_sub_0_o[2]~14 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_25_sub_0_o[1]~13 ),
	.combout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[2]~14_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[2]~15 ));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[2]~14 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[2]~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_25_sub_0_o[3]~16 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_25_sub_0_o[2]~15 ),
	.combout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[3]~16_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[3]~17 ));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[3]~16 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[3]~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_25_sub_0_o[4]~18 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_25_sub_0_o[3]~17 ),
	.combout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[4]~18_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[4]~19 ));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[4]~18 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[4]~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_25_sub_0_o[5]~20 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_25_sub_0_o[4]~19 ),
	.combout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[5]~20_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[5]~21 ));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[5]~20 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[5]~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_25_sub_0_o[6]~22 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_25_sub_0_o[5]~21 ),
	.combout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[6]~22_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[6]~23 ));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[6]~22 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[6]~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_25_sub_0_o[7]~24 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_25_sub_0_o[6]~23 ),
	.combout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[7]~24_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[7]~25 ));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[7]~24 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[7]~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_25_sub_0_o[8]~26 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_25_sub_0_o[7]~25 ),
	.combout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[8]~26_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[8]~27 ));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[8]~26 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[8]~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_25_sub_0_o[9]~28 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_25_sub_0_o[8]~27 ),
	.combout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[9]~28_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[9]~29 ));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[9]~28 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[9]~28 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_25_sub_0_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_25_sub_0_o[9]~28_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_25_sub_0_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_25_sub_0_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_25_sub_0_o[8]~26_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_25_sub_0_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_25_sub_0_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_25_sub_0_o[7]~24_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_25_sub_0_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_25_sub_0_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_25_sub_0_o[6]~22_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_25_sub_0_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_25_sub_0_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_25_sub_0_o[5]~20_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_25_sub_0_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_25_sub_0_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_25_sub_0_o[4]~18_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_25_sub_0_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_25_sub_0_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_25_sub_0_o[3]~16_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_25_sub_0_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_25_sub_0_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_25_sub_0_o[2]~14_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_25_sub_0_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_25_sub_0_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_25_sub_0_o[1]~12_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_25_sub_0_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_25_sub_0_o[0] (
	.clk(clk),
	.d(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_25_sub_0_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_12_o[0]~14 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][0]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_25_sub_0_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_add0_12_o[0]~14_combout ),
	.cout(\u0_m0_wo0_mtree_add0_12_o[0]~15 ));
defparam \u0_m0_wo0_mtree_add0_12_o[0]~14 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_add0_12_o[0]~14 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_12_o[1]~16 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][1]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_25_sub_0_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_12_o[0]~15 ),
	.combout(\u0_m0_wo0_mtree_add0_12_o[1]~16_combout ),
	.cout(\u0_m0_wo0_mtree_add0_12_o[1]~17 ));
defparam \u0_m0_wo0_mtree_add0_12_o[1]~16 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_12_o[1]~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_12_o[2]~18 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][2]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_25_sub_0_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_12_o[1]~17 ),
	.combout(\u0_m0_wo0_mtree_add0_12_o[2]~18_combout ),
	.cout(\u0_m0_wo0_mtree_add0_12_o[2]~19 ));
defparam \u0_m0_wo0_mtree_add0_12_o[2]~18 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_12_o[2]~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_12_o[3]~20 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][3]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_25_sub_0_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_12_o[2]~19 ),
	.combout(\u0_m0_wo0_mtree_add0_12_o[3]~20_combout ),
	.cout(\u0_m0_wo0_mtree_add0_12_o[3]~21 ));
defparam \u0_m0_wo0_mtree_add0_12_o[3]~20 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_12_o[3]~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_12_o[4]~22 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][4]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_25_sub_0_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_12_o[3]~21 ),
	.combout(\u0_m0_wo0_mtree_add0_12_o[4]~22_combout ),
	.cout(\u0_m0_wo0_mtree_add0_12_o[4]~23 ));
defparam \u0_m0_wo0_mtree_add0_12_o[4]~22 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_12_o[4]~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_12_o[5]~24 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][5]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_25_sub_0_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_12_o[4]~23 ),
	.combout(\u0_m0_wo0_mtree_add0_12_o[5]~24_combout ),
	.cout(\u0_m0_wo0_mtree_add0_12_o[5]~25 ));
defparam \u0_m0_wo0_mtree_add0_12_o[5]~24 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_12_o[5]~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_12_o[6]~26 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][6]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_25_sub_0_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_12_o[5]~25 ),
	.combout(\u0_m0_wo0_mtree_add0_12_o[6]~26_combout ),
	.cout(\u0_m0_wo0_mtree_add0_12_o[6]~27 ));
defparam \u0_m0_wo0_mtree_add0_12_o[6]~26 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_12_o[6]~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_12_o[7]~28 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][7]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_25_sub_0_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_12_o[6]~27 ),
	.combout(\u0_m0_wo0_mtree_add0_12_o[7]~28_combout ),
	.cout(\u0_m0_wo0_mtree_add0_12_o[7]~29 ));
defparam \u0_m0_wo0_mtree_add0_12_o[7]~28 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_12_o[7]~28 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_12_o[8]~30 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][8]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_25_sub_0_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_12_o[7]~29 ),
	.combout(\u0_m0_wo0_mtree_add0_12_o[8]~30_combout ),
	.cout(\u0_m0_wo0_mtree_add0_12_o[8]~31 ));
defparam \u0_m0_wo0_mtree_add0_12_o[8]~30 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_12_o[8]~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_12_o[9]~32 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][9]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_25_sub_0_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_12_o[8]~31 ),
	.combout(\u0_m0_wo0_mtree_add0_12_o[9]~32_combout ),
	.cout(\u0_m0_wo0_mtree_add0_12_o[9]~33 ));
defparam \u0_m0_wo0_mtree_add0_12_o[9]~32 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_12_o[9]~32 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add0_12_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_12_o[9]~32_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_12_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_12_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_12_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_2_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[8]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_12_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_12_o[8]~30_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_12_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_12_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_12_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_2_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[7]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_12_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_12_o[7]~28_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_12_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_12_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_12_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_2_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[6]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_12_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_12_o[6]~26_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_12_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_12_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_12_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_2_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[5]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_12_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_12_o[5]~24_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_12_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_12_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_12_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_2_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[4]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_12_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_12_o[4]~22_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_12_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_12_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_12_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_2_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[3]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_12_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_12_o[3]~20_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_12_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_12_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_12_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_2_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[2]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_12_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_12_o[2]~18_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_12_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_12_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_12_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_2_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[1]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_12_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_12_o[1]~16_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_12_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_12_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_12_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_2_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[0]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_12_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_12_o[0]~14_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_12_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_12_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_12_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[0]~21 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\u0_m0_wo0_mtree_add3_1_o[0]~21_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[0]~22 ));
defparam \u0_m0_wo0_mtree_add3_1_o[0]~21 .lut_mask = 16'h6688;
defparam \u0_m0_wo0_mtree_add3_1_o[0]~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[1]~23 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[1]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_1_o[0]~22 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[1]~23_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[1]~24 ));
defparam \u0_m0_wo0_mtree_add3_1_o[1]~23 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_1_o[1]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[2]~25 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[2]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_1_o[1]~24 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[2]~25_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[2]~26 ));
defparam \u0_m0_wo0_mtree_add3_1_o[2]~25 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add3_1_o[2]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[3]~27 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[3]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_1_o[2]~26 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[3]~27_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[3]~28 ));
defparam \u0_m0_wo0_mtree_add3_1_o[3]~27 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_1_o[3]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[4]~29 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[4]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_1_o[3]~28 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[4]~29_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[4]~30 ));
defparam \u0_m0_wo0_mtree_add3_1_o[4]~29 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add3_1_o[4]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[5]~31 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[5]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_1_o[4]~30 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[5]~31_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[5]~32 ));
defparam \u0_m0_wo0_mtree_add3_1_o[5]~31 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_1_o[5]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[6]~33 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[6]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_1_o[5]~32 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[6]~33_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[6]~34 ));
defparam \u0_m0_wo0_mtree_add3_1_o[6]~33 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add3_1_o[6]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[7]~35 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[7]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_1_o[6]~34 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[7]~35_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[7]~36 ));
defparam \u0_m0_wo0_mtree_add3_1_o[7]~35 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_1_o[7]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[8]~37 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[8]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_1_o[7]~36 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[8]~37_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[8]~38 ));
defparam \u0_m0_wo0_mtree_add3_1_o[8]~37 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add3_1_o[8]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[9]~39 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[9]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_1_o[8]~38 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[9]~39_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[9]~40 ));
defparam \u0_m0_wo0_mtree_add3_1_o[9]~39 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_1_o[9]~39 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add3_1_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[9]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[9] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_0_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[8]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_1_o[8] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[8]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[8]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[8] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[8] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_0_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[7]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_1_o[7] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[7]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[7]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[7] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[7] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_0_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[6]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_1_o[6] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[6]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[6]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[6] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[6] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_0_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[5]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_1_o[5] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[5]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[5]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[5] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[5] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_0_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[4]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_1_o[4] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[4]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[4]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[4] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[4] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_0_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[3]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_1_o[3] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[3]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[3]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[3] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[3] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_0_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[2]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_1_o[2] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[2]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[2]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[2] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[2] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_0_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[1]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_1_o[1] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[1]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[1]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[1] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[1] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_0_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[0]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[0] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_1_o[0] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[0]~21_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[0]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[0] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[0] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[9]~13 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[0]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\u0_m0_wo0_mtree_add4_0_o[9]~13_cout ));
defparam \u0_m0_wo0_mtree_add4_0_o[9]~13 .lut_mask = 16'h0088;
defparam \u0_m0_wo0_mtree_add4_0_o[9]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[9]~15 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[1]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add4_0_o[9]~13_cout ),
	.combout(),
	.cout(\u0_m0_wo0_mtree_add4_0_o[9]~15_cout ));
defparam \u0_m0_wo0_mtree_add4_0_o[9]~15 .lut_mask = 16'h0017;
defparam \u0_m0_wo0_mtree_add4_0_o[9]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[9]~17 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[2]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add4_0_o[9]~15_cout ),
	.combout(),
	.cout(\u0_m0_wo0_mtree_add4_0_o[9]~17_cout ));
defparam \u0_m0_wo0_mtree_add4_0_o[9]~17 .lut_mask = 16'h008E;
defparam \u0_m0_wo0_mtree_add4_0_o[9]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[9]~19 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[3]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add4_0_o[9]~17_cout ),
	.combout(),
	.cout(\u0_m0_wo0_mtree_add4_0_o[9]~19_cout ));
defparam \u0_m0_wo0_mtree_add4_0_o[9]~19 .lut_mask = 16'h0017;
defparam \u0_m0_wo0_mtree_add4_0_o[9]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[9]~21 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[4]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add4_0_o[9]~19_cout ),
	.combout(),
	.cout(\u0_m0_wo0_mtree_add4_0_o[9]~21_cout ));
defparam \u0_m0_wo0_mtree_add4_0_o[9]~21 .lut_mask = 16'h008E;
defparam \u0_m0_wo0_mtree_add4_0_o[9]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[9]~23 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[5]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add4_0_o[9]~21_cout ),
	.combout(),
	.cout(\u0_m0_wo0_mtree_add4_0_o[9]~23_cout ));
defparam \u0_m0_wo0_mtree_add4_0_o[9]~23 .lut_mask = 16'h0017;
defparam \u0_m0_wo0_mtree_add4_0_o[9]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[9]~25 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[6]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add4_0_o[9]~23_cout ),
	.combout(),
	.cout(\u0_m0_wo0_mtree_add4_0_o[9]~25_cout ));
defparam \u0_m0_wo0_mtree_add4_0_o[9]~25 .lut_mask = 16'h008E;
defparam \u0_m0_wo0_mtree_add4_0_o[9]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[9]~27 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[7]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add4_0_o[9]~25_cout ),
	.combout(),
	.cout(\u0_m0_wo0_mtree_add4_0_o[9]~27_cout ));
defparam \u0_m0_wo0_mtree_add4_0_o[9]~27 .lut_mask = 16'h0017;
defparam \u0_m0_wo0_mtree_add4_0_o[9]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[9]~29 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[8]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add4_0_o[9]~27_cout ),
	.combout(),
	.cout(\u0_m0_wo0_mtree_add4_0_o[9]~29_cout ));
defparam \u0_m0_wo0_mtree_add4_0_o[9]~29 .lut_mask = 16'h008E;
defparam \u0_m0_wo0_mtree_add4_0_o[9]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[9]~30 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[9]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add4_0_o[9]~29_cout ),
	.combout(\u0_m0_wo0_mtree_add4_0_o[9]~30_combout ),
	.cout(\u0_m0_wo0_mtree_add4_0_o[9]~31 ));
defparam \u0_m0_wo0_mtree_add4_0_o[9]~30 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add4_0_o[9]~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_5_sub_0_o[10]~30 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_5_sub_0_o[9]~29 ),
	.combout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[10]~30_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[10]~31 ));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[10]~30 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[10]~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_5_sub_0_o[11]~32 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_5_sub_0_o[10]~31 ),
	.combout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[11]~32_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[11]~33 ));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[11]~32 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[11]~32 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_5_sub_0_o[12]~34 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr25|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_5_sub_0_o[11]~33 ),
	.combout(\u0_m0_wo0_mtree_mult1_5_sub_0_o[12]~34_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[12]~34 .lut_mask = 16'hA5A5;
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[12]~34 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_5_sub_0_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_5_sub_0_o[12]~34_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_5_sub_0_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_5_sub_0_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_5_sub_0_o[11]~32_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_5_sub_0_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_5_sub_0_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_5_sub_0_o[10]~30_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_5_sub_0_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_5_sub_0_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_1_o[10]~34 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][10]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_5_sub_0_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_1_o[9]~33 ),
	.combout(\u0_m0_wo0_mtree_add1_1_o[10]~34_combout ),
	.cout(\u0_m0_wo0_mtree_add1_1_o[10]~35 ));
defparam \u0_m0_wo0_mtree_add1_1_o[10]~34 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_1_o[10]~34 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_1_o[11]~36 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_5_sub_0_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_1_o[10]~35 ),
	.combout(\u0_m0_wo0_mtree_add1_1_o[11]~36_combout ),
	.cout(\u0_m0_wo0_mtree_add1_1_o[11]~37 ));
defparam \u0_m0_wo0_mtree_add1_1_o[11]~36 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_1_o[11]~36 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_1_o[12]~38 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_5_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_1_o[11]~37 ),
	.combout(\u0_m0_wo0_mtree_add1_1_o[12]~38_combout ),
	.cout(\u0_m0_wo0_mtree_add1_1_o[12]~39 ));
defparam \u0_m0_wo0_mtree_add1_1_o[12]~38 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_1_o[12]~38 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_1_o[15]~40 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_5_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_add1_1_o[12]~39 ),
	.combout(\u0_m0_wo0_mtree_add1_1_o[15]~40_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_add1_1_o[15]~40 .lut_mask = 16'h9696;
defparam \u0_m0_wo0_mtree_add1_1_o[15]~40 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add1_1_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_1_o[15]~40_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_1_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_1_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_1_o[15] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_8_sub_1_o[10]~29 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][8]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_8_sub_1_o[9]~28 ),
	.combout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[10]~29_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[10]~30 ));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[10]~29 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[10]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_8_sub_1_o[11]~31 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][9]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_8_sub_1_o[10]~30 ),
	.combout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[11]~31_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[11]~32 ));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[11]~31 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[11]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_8_sub_1_o[12]~33 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][10]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr22|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_8_sub_1_o[11]~32 ),
	.combout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[12]~33_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[12]~34 ));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[12]~33 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[12]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_8_sub_1_o[13]~35 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_8_sub_1_o[12]~34 ),
	.combout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[13]~35_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[13]~36 ));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[13]~35 .lut_mask = 16'h0F0F;
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[13]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_8_sub_1_o[14]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_8_sub_1_o[13]~36 ),
	.combout(\u0_m0_wo0_mtree_mult1_8_sub_1_o[14]~37_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[14]~37 .lut_mask = 16'hF0F0;
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[14]~37 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_8_sub_1_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_8_sub_1_o[14]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_8_sub_1_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[14] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_9_add_1_o[9]~29 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][8]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_9_add_1_o[8]~28 ),
	.combout(\u0_m0_wo0_mtree_mult1_9_add_1_o[9]~29_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_9_add_1_o[9]~30 ));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[9]~29 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[9]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_9_add_1_o[10]~31 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][10]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_9_add_1_o[9]~30 ),
	.combout(\u0_m0_wo0_mtree_mult1_9_add_1_o[10]~31_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_9_add_1_o[10]~32 ));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[10]~31 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[10]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_9_add_1_o[11]~33 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][10]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_9_add_1_o[10]~32 ),
	.combout(\u0_m0_wo0_mtree_mult1_9_add_1_o[11]~33_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_9_add_1_o[11]~34 ));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[11]~33 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[11]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_9_add_1_o[12]~35 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr21|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_9_add_1_o[11]~34 ),
	.combout(\u0_m0_wo0_mtree_mult1_9_add_1_o[12]~35_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_9_add_1_o[12]~36 ));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[12]~35 .lut_mask = 16'hF0AA;
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[12]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_9_add_1_o[13]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_9_add_1_o[12]~36 ),
	.combout(\u0_m0_wo0_mtree_mult1_9_add_1_o[13]~37_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[13]~37 .lut_mask = 16'hF0F0;
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[13]~37 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_9_add_1_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_9_add_1_o[13]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_9_add_1_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_8_sub_1_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_8_sub_1_o[13]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_8_sub_1_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_9_add_1_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_9_add_1_o[12]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_9_add_1_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_8_sub_1_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_8_sub_1_o[12]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_8_sub_1_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_9_add_1_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_9_add_1_o[11]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_9_add_1_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_8_sub_1_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_8_sub_1_o[11]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_8_sub_1_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_9_add_1_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_9_add_1_o[10]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_9_add_1_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[10] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_8_sub_1_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_8_sub_1_o[10]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_8_sub_1_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_8_sub_1_o[10] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_9_add_1_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_9_add_1_o[9]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_9_add_1_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_9_add_1_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_4_o[10]~33 (
	.dataa(\u0_m0_wo0_mtree_mult1_8_sub_1_o[10]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_9_add_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_4_o[9]~32 ),
	.combout(\u0_m0_wo0_mtree_add0_4_o[10]~33_combout ),
	.cout(\u0_m0_wo0_mtree_add0_4_o[10]~34 ));
defparam \u0_m0_wo0_mtree_add0_4_o[10]~33 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_4_o[10]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_4_o[11]~35 (
	.dataa(\u0_m0_wo0_mtree_mult1_8_sub_1_o[11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_9_add_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_4_o[10]~34 ),
	.combout(\u0_m0_wo0_mtree_add0_4_o[11]~35_combout ),
	.cout(\u0_m0_wo0_mtree_add0_4_o[11]~36 ));
defparam \u0_m0_wo0_mtree_add0_4_o[11]~35 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_4_o[11]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_4_o[12]~37 (
	.dataa(\u0_m0_wo0_mtree_mult1_8_sub_1_o[12]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_9_add_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_4_o[11]~36 ),
	.combout(\u0_m0_wo0_mtree_add0_4_o[12]~37_combout ),
	.cout(\u0_m0_wo0_mtree_add0_4_o[12]~38 ));
defparam \u0_m0_wo0_mtree_add0_4_o[12]~37 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_4_o[12]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_4_o[13]~39 (
	.dataa(\u0_m0_wo0_mtree_mult1_8_sub_1_o[13]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_9_add_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_4_o[12]~38 ),
	.combout(\u0_m0_wo0_mtree_add0_4_o[13]~39_combout ),
	.cout(\u0_m0_wo0_mtree_add0_4_o[13]~40 ));
defparam \u0_m0_wo0_mtree_add0_4_o[13]~39 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_4_o[13]~39 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_4_o[14]~41 (
	.dataa(\u0_m0_wo0_mtree_mult1_8_sub_1_o[14]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_9_add_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_4_o[13]~40 ),
	.combout(\u0_m0_wo0_mtree_add0_4_o[14]~41_combout ),
	.cout(\u0_m0_wo0_mtree_add0_4_o[14]~42 ));
defparam \u0_m0_wo0_mtree_add0_4_o[14]~41 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_4_o[14]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_4_o[15]~43 (
	.dataa(\u0_m0_wo0_mtree_mult1_8_sub_1_o[14]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_9_add_1_o[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_add0_4_o[14]~42 ),
	.combout(\u0_m0_wo0_mtree_add0_4_o[15]~43_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_add0_4_o[15]~43 .lut_mask = 16'h6969;
defparam \u0_m0_wo0_mtree_add0_4_o[15]~43 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add0_4_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_4_o[15]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_4_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_4_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_4_o[15] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_0_o[10]~30 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_0_o[9]~29 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[10]~30_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[10]~31 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[10]~30 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[10]~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_0_o[11]~32 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_0_o[10]~31 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[11]~32_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[11]~33 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[11]~32 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[11]~32 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_0_o[12]~34 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr20|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_0_o[11]~33 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_0_o[12]~34_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[12]~34 .lut_mask = 16'hA5A5;
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[12]~34 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_0_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_0_o[12]~34_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_0_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_0_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_0_o[11]~32_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_0_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_0_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_0_o[10]~30_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_0_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_0_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_2_o[10]~29 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][8]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_0_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_2_o[9]~28 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[10]~29_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[10]~30 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[10]~29 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[10]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_2_o[11]~31 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][9]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_0_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_2_o[10]~30 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[11]~31_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[11]~32 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[11]~31 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[11]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_2_o[12]~33 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][10]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_2_o[11]~32 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[12]~33_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[12]~34 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[12]~33 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[12]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_2_o[13]~35 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_2_o[12]~34 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[13]~35_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[13]~36 ));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[13]~35 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[13]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_10_sub_2_o[14]~37 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_10_sub_2_o[13]~36 ),
	.combout(\u0_m0_wo0_mtree_mult1_10_sub_2_o[14]~37_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[14]~37 .lut_mask = 16'h9696;
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[14]~37 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_2_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_2_o[14]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_2_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_4_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_4_o[14]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_4_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_4_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_4_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_4_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_4_o[13]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_4_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_4_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_4_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_2_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_2_o[13]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_2_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_4_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_4_o[12]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_4_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_4_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_4_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_2_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_2_o[12]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_2_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_4_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_4_o[11]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_4_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_4_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_4_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_2_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_2_o[11]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_2_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_4_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_4_o[10]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_4_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_4_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_4_o[10] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_10_sub_2_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_10_sub_2_o[10]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_10_sub_2_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_10_sub_2_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_2_o[10]~37 (
	.dataa(\u0_m0_wo0_mtree_add0_4_o[10]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_2_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_2_o[9]~36 ),
	.combout(\u0_m0_wo0_mtree_add1_2_o[10]~37_combout ),
	.cout(\u0_m0_wo0_mtree_add1_2_o[10]~38 ));
defparam \u0_m0_wo0_mtree_add1_2_o[10]~37 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_2_o[10]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_2_o[11]~39 (
	.dataa(\u0_m0_wo0_mtree_add0_4_o[11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_2_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_2_o[10]~38 ),
	.combout(\u0_m0_wo0_mtree_add1_2_o[11]~39_combout ),
	.cout(\u0_m0_wo0_mtree_add1_2_o[11]~40 ));
defparam \u0_m0_wo0_mtree_add1_2_o[11]~39 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_2_o[11]~39 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_2_o[12]~41 (
	.dataa(\u0_m0_wo0_mtree_add0_4_o[12]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_2_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_2_o[11]~40 ),
	.combout(\u0_m0_wo0_mtree_add1_2_o[12]~41_combout ),
	.cout(\u0_m0_wo0_mtree_add1_2_o[12]~42 ));
defparam \u0_m0_wo0_mtree_add1_2_o[12]~41 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_2_o[12]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_2_o[13]~43 (
	.dataa(\u0_m0_wo0_mtree_add0_4_o[13]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_2_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_2_o[12]~42 ),
	.combout(\u0_m0_wo0_mtree_add1_2_o[13]~43_combout ),
	.cout(\u0_m0_wo0_mtree_add1_2_o[13]~44 ));
defparam \u0_m0_wo0_mtree_add1_2_o[13]~43 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_2_o[13]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_2_o[14]~45 (
	.dataa(\u0_m0_wo0_mtree_add0_4_o[14]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_2_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_2_o[13]~44 ),
	.combout(\u0_m0_wo0_mtree_add1_2_o[14]~45_combout ),
	.cout(\u0_m0_wo0_mtree_add1_2_o[14]~46 ));
defparam \u0_m0_wo0_mtree_add1_2_o[14]~45 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_2_o[14]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_2_o[15]~47 (
	.dataa(\u0_m0_wo0_mtree_add0_4_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_2_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_2_o[14]~46 ),
	.combout(\u0_m0_wo0_mtree_add1_2_o[15]~47_combout ),
	.cout(\u0_m0_wo0_mtree_add1_2_o[15]~48 ));
defparam \u0_m0_wo0_mtree_add1_2_o[15]~47 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_2_o[15]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_2_o[17]~49 (
	.dataa(\u0_m0_wo0_mtree_add0_4_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_10_sub_2_o[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_add1_2_o[15]~48 ),
	.combout(\u0_m0_wo0_mtree_add1_2_o[17]~49_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_add1_2_o[17]~49 .lut_mask = 16'h6969;
defparam \u0_m0_wo0_mtree_add1_2_o[17]~49 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add1_2_o[17] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_2_o[17]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_2_o[17]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_2_o[17] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_2_o[17] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_1_o[10]~31 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][10]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_1_o[9]~30 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_1_o[10]~31_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_1_o[10]~32 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[10]~31 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[10]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_1_o[11]~33 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][10]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_1_o[10]~32 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_1_o[11]~33_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_1_o[11]~34 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[11]~33 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[11]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_1_o[12]~35 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr18|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_1_o[11]~34 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_1_o[12]~35_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_1_o[12]~36 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[12]~35 .lut_mask = 16'hF0AA;
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[12]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_1_o[13]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_1_o[12]~36 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_1_o[13]~37_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[13]~37 .lut_mask = 16'hF0F0;
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[13]~37 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_12_add_1_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_1_o[13]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_1_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_1_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_1_o[12]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_1_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_1_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_1_o[11]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_1_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_1_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_1_o[10]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_1_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_3_o[10]~27 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][7]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_12_add_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_3_o[9]~26 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_3_o[10]~27_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_3_o[10]~28 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[10]~27 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[10]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_3_o[11]~29 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][8]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_12_add_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_3_o[10]~28 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_3_o[11]~29_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_3_o[11]~30 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[11]~29 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[11]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_3_o[12]~31 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][9]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_12_add_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_3_o[11]~30 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_3_o[12]~31_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_3_o[12]~32 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[12]~31 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[12]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_3_o[13]~33 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][10]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_12_add_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_3_o[12]~32 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_3_o[13]~33_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_3_o[13]~34 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[13]~33 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[13]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_3_o[14]~35 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_12_add_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_3_o[13]~34 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_3_o[14]~35_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_12_add_3_o[14]~36 ));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[14]~35 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[14]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_12_add_3_o[15]~37 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_12_add_1_o[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_12_add_3_o[14]~36 ),
	.combout(\u0_m0_wo0_mtree_mult1_12_add_3_o[15]~37_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[15]~37 .lut_mask = 16'h6969;
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[15]~37 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_12_add_3_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_3_o[15]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_3_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[15] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_1_o[10]~33 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][7]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_1_o[9]~32 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[10]~33_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[10]~34 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[10]~33 .lut_mask = 16'h694D;
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[10]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_1_o[11]~35 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][8]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_1_o[10]~34 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[11]~35_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[11]~36 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[11]~35 .lut_mask = 16'h962B;
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[11]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_1_o[12]~37 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][9]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_1_o[11]~36 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[12]~37_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[12]~38 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[12]~37 .lut_mask = 16'h694D;
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[12]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_1_o[13]~39 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][10]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr17|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_1_o[12]~38 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[13]~39_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[13]~40 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[13]~39 .lut_mask = 16'h962B;
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[13]~39 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_1_o[14]~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_1_o[13]~40 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[14]~41_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[14]~42 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[14]~41 .lut_mask = 16'h0F0F;
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[14]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_1_o[15]~43 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_1_o[14]~42 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_1_o[15]~43_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[15]~43 .lut_mask = 16'hF0F0;
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[15]~43 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_1_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[15]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_1_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_1_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[14]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_1_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_1_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[13]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_1_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_1_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[12]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_1_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_1_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[11]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_1_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_1_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_1_o[10]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_1_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_3_o[10]~23 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][5]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_3_o[9]~22 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[10]~23_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[10]~24 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[10]~23 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[10]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_3_o[11]~25 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][6]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_3_o[10]~24 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[11]~25_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[11]~26 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[11]~25 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[11]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_3_o[12]~27 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][7]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_3_o[11]~26 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[12]~27_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[12]~28 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[12]~27 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[12]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_3_o[13]~29 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][8]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_3_o[12]~28 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[13]~29_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[13]~30 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[13]~29 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[13]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_3_o[14]~31 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][9]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_3_o[13]~30 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[14]~31_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[14]~32 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[14]~31 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[14]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_3_o[15]~33 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][10]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_1_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_3_o[14]~32 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[15]~33_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[15]~34 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[15]~33 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[15]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_3_o[16]~35 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_1_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_3_o[15]~34 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[16]~35_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[16]~36 ));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[16]~35 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[16]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_13_sub_3_o[17]~37 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_1_o[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_13_sub_3_o[16]~36 ),
	.combout(\u0_m0_wo0_mtree_mult1_13_sub_3_o[17]~37_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[17]~37 .lut_mask = 16'h9696;
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[17]~37 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_3_o[17] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_3_o[17]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_3_o[17]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[17] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[17] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_3_o[16] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_3_o[16]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_3_o[16]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[16] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[16] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_3_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_3_o[15]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_3_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_3_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_3_o[14]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_3_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_3_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_3_o[14]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_3_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_3_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_3_o[13]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_3_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_3_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_3_o[13]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_3_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_3_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_3_o[12]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_3_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_3_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_3_o[12]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_3_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_3_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_3_o[11]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_3_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_3_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_3_o[11]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_3_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_12_add_3_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_12_add_3_o[10]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_12_add_3_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_12_add_3_o[10] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_13_sub_3_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_13_sub_3_o[10]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_13_sub_3_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_13_sub_3_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_6_o[10]~39 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_3_o[10]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_3_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_6_o[9]~38 ),
	.combout(\u0_m0_wo0_mtree_add0_6_o[10]~39_combout ),
	.cout(\u0_m0_wo0_mtree_add0_6_o[10]~40 ));
defparam \u0_m0_wo0_mtree_add0_6_o[10]~39 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_6_o[10]~39 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_6_o[11]~41 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_3_o[11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_3_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_6_o[10]~40 ),
	.combout(\u0_m0_wo0_mtree_add0_6_o[11]~41_combout ),
	.cout(\u0_m0_wo0_mtree_add0_6_o[11]~42 ));
defparam \u0_m0_wo0_mtree_add0_6_o[11]~41 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_6_o[11]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_6_o[12]~43 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_3_o[12]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_3_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_6_o[11]~42 ),
	.combout(\u0_m0_wo0_mtree_add0_6_o[12]~43_combout ),
	.cout(\u0_m0_wo0_mtree_add0_6_o[12]~44 ));
defparam \u0_m0_wo0_mtree_add0_6_o[12]~43 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_6_o[12]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_6_o[13]~45 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_3_o[13]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_3_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_6_o[12]~44 ),
	.combout(\u0_m0_wo0_mtree_add0_6_o[13]~45_combout ),
	.cout(\u0_m0_wo0_mtree_add0_6_o[13]~46 ));
defparam \u0_m0_wo0_mtree_add0_6_o[13]~45 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_6_o[13]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_6_o[14]~47 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_3_o[14]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_3_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_6_o[13]~46 ),
	.combout(\u0_m0_wo0_mtree_add0_6_o[14]~47_combout ),
	.cout(\u0_m0_wo0_mtree_add0_6_o[14]~48 ));
defparam \u0_m0_wo0_mtree_add0_6_o[14]~47 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_6_o[14]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_6_o[15]~49 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_3_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_3_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_6_o[14]~48 ),
	.combout(\u0_m0_wo0_mtree_add0_6_o[15]~49_combout ),
	.cout(\u0_m0_wo0_mtree_add0_6_o[15]~50 ));
defparam \u0_m0_wo0_mtree_add0_6_o[15]~49 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_6_o[15]~49 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_6_o[16]~51 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_3_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_3_o[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_6_o[15]~50 ),
	.combout(\u0_m0_wo0_mtree_add0_6_o[16]~51_combout ),
	.cout(\u0_m0_wo0_mtree_add0_6_o[16]~52 ));
defparam \u0_m0_wo0_mtree_add0_6_o[16]~51 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_6_o[16]~51 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_6_o[17]~53 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_3_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_3_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_6_o[16]~52 ),
	.combout(\u0_m0_wo0_mtree_add0_6_o[17]~53_combout ),
	.cout(\u0_m0_wo0_mtree_add0_6_o[17]~54 ));
defparam \u0_m0_wo0_mtree_add0_6_o[17]~53 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_6_o[17]~53 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_6_o[18]~55 (
	.dataa(\u0_m0_wo0_mtree_mult1_12_add_3_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_13_sub_3_o[17]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_add0_6_o[17]~54 ),
	.combout(\u0_m0_wo0_mtree_add0_6_o[18]~55_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_add0_6_o[18]~55 .lut_mask = 16'h6969;
defparam \u0_m0_wo0_mtree_add0_6_o[18]~55 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add0_6_o[18] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_6_o[18]~55_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_6_o[18]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_6_o[18] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_6_o[18] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_1_o[10]~29 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][8]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_1_o[9]~28 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_1_o[10]~29_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_1_o[10]~30 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[10]~29 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[10]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_1_o[11]~31 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][9]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_1_o[10]~30 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_1_o[11]~31_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_1_o[11]~32 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[11]~31 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[11]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_1_o[12]~33 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][10]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_1_o[11]~32 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_1_o[12]~33_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_1_o[12]~34 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[12]~33 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[12]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_1_o[13]~35 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr16|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_1_o[12]~34 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_1_o[13]~35_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_1_o[13]~36 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[13]~35 .lut_mask = 16'hF0AA;
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[13]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_1_o[14]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_1_o[13]~36 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_1_o[14]~37_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[14]~37 .lut_mask = 16'hF0F0;
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[14]~37 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_14_add_1_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_1_o[14]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_1_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_1_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_1_o[13]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_1_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_1_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_1_o[12]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_1_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_1_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_1_o[11]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_1_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_1_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_1_o[10]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_1_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_3_o[10]~23 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][5]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_14_add_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_3_o[9]~22 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_3_o[10]~23_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_3_o[10]~24 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[10]~23 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[10]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_3_o[11]~25 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][6]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_14_add_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_3_o[10]~24 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_3_o[11]~25_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_3_o[11]~26 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[11]~25 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[11]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_3_o[12]~27 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][7]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_14_add_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_3_o[11]~26 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_3_o[12]~27_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_3_o[12]~28 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[12]~27 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[12]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_3_o[13]~29 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][8]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_14_add_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_3_o[12]~28 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_3_o[13]~29_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_3_o[13]~30 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[13]~29 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[13]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_3_o[14]~31 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][9]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_14_add_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_3_o[13]~30 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_3_o[14]~31_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_3_o[14]~32 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[14]~31 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[14]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_3_o[15]~33 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][10]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_14_add_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_3_o[14]~32 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_3_o[15]~33_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_3_o[15]~34 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[15]~33 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[15]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_3_o[16]~35 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_14_add_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_3_o[15]~34 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_3_o[16]~35_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_14_add_3_o[16]~36 ));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[16]~35 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[16]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_14_add_3_o[17]~37 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_14_add_1_o[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_14_add_3_o[16]~36 ),
	.combout(\u0_m0_wo0_mtree_mult1_14_add_3_o[17]~37_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[17]~37 .lut_mask = 16'h6969;
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[17]~37 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_14_add_3_o[17] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_3_o[17]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_3_o[17]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[17] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[17] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_15_sub_1_o[10]~37 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][3]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_15_sub_1_o[9]~36 ),
	.combout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[10]~37_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[10]~38 ));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[10]~37 .lut_mask = 16'h694D;
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[10]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_15_sub_1_o[11]~39 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][4]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_15_sub_1_o[10]~38 ),
	.combout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[11]~39_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[11]~40 ));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[11]~39 .lut_mask = 16'h962B;
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[11]~39 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_15_sub_1_o[12]~41 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][5]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_15_sub_1_o[11]~40 ),
	.combout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[12]~41_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[12]~42 ));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[12]~41 .lut_mask = 16'h694D;
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[12]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_15_sub_1_o[13]~43 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][6]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_15_sub_1_o[12]~42 ),
	.combout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[13]~43_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[13]~44 ));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[13]~43 .lut_mask = 16'h962B;
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[13]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_15_sub_1_o[14]~45 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][7]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_15_sub_1_o[13]~44 ),
	.combout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[14]~45_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[14]~46 ));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[14]~45 .lut_mask = 16'h694D;
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[14]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_15_sub_1_o[15]~47 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][8]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_15_sub_1_o[14]~46 ),
	.combout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[15]~47_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[15]~48 ));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[15]~47 .lut_mask = 16'h962B;
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[15]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_15_sub_1_o[16]~49 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][9]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_15_sub_1_o[15]~48 ),
	.combout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[16]~49_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[16]~50 ));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[16]~49 .lut_mask = 16'h694D;
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[16]~49 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_15_sub_1_o[17]~51 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][10]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_15_sub_1_o[16]~50 ),
	.combout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[17]~51_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[17]~52 ));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[17]~51 .lut_mask = 16'h962B;
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[17]~51 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_15_sub_1_o[18]~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_15_sub_1_o[17]~52 ),
	.combout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[18]~53_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[18]~54 ));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[18]~53 .lut_mask = 16'h0F0F;
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[18]~53 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_15_sub_1_o[19]~55 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_15_sub_1_o[18]~54 ),
	.combout(\u0_m0_wo0_mtree_mult1_15_sub_1_o[19]~55_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[19]~55 .lut_mask = 16'hF0F0;
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[19]~55 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[19] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_15_sub_1_o[19]~55_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[19]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[19] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[19] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[18] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_15_sub_1_o[18]~53_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[18]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[18] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[18] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[17] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_15_sub_1_o[17]~51_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[17]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[17] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[17] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_3_o[16] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_3_o[16]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_3_o[16]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[16] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[16] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[16] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_15_sub_1_o[16]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[16]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[16] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[16] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_3_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_3_o[15]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_3_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_15_sub_1_o[15]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_3_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_3_o[14]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_3_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_15_sub_1_o[14]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_3_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_3_o[13]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_3_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_15_sub_1_o[13]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_3_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_3_o[12]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_3_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_15_sub_1_o[12]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_3_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_3_o[11]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_3_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_15_sub_1_o[11]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_14_add_3_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_14_add_3_o[10]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_14_add_3_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_14_add_3_o[10] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_15_sub_1_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_15_sub_1_o[10]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_15_sub_1_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_15_sub_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[10]~41 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[10]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_7_o[9]~40 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[10]~41_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[10]~42 ));
defparam \u0_m0_wo0_mtree_add0_7_o[10]~41 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_7_o[10]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[11]~43 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_7_o[10]~42 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[11]~43_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[11]~44 ));
defparam \u0_m0_wo0_mtree_add0_7_o[11]~43 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_7_o[11]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[12]~45 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[12]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_7_o[11]~44 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[12]~45_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[12]~46 ));
defparam \u0_m0_wo0_mtree_add0_7_o[12]~45 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_7_o[12]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[13]~47 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[13]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_7_o[12]~46 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[13]~47_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[13]~48 ));
defparam \u0_m0_wo0_mtree_add0_7_o[13]~47 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_7_o[13]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[14]~49 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[14]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_7_o[13]~48 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[14]~49_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[14]~50 ));
defparam \u0_m0_wo0_mtree_add0_7_o[14]~49 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_7_o[14]~49 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[15]~51 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_7_o[14]~50 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[15]~51_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[15]~52 ));
defparam \u0_m0_wo0_mtree_add0_7_o[15]~51 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_7_o[15]~51 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[16]~53 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[16]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_7_o[15]~52 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[16]~53_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[16]~54 ));
defparam \u0_m0_wo0_mtree_add0_7_o[16]~53 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_7_o[16]~53 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[17]~55 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[17]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_7_o[16]~54 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[17]~55_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[17]~56 ));
defparam \u0_m0_wo0_mtree_add0_7_o[17]~55 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_7_o[17]~55 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[18]~57 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[17]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[18]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_7_o[17]~56 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[18]~57_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[18]~58 ));
defparam \u0_m0_wo0_mtree_add0_7_o[18]~57 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_7_o[18]~57 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[19]~59 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[17]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[19]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_7_o[18]~58 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[19]~59_combout ),
	.cout(\u0_m0_wo0_mtree_add0_7_o[19]~60 ));
defparam \u0_m0_wo0_mtree_add0_7_o[19]~59 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_7_o[19]~59 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_7_o[20]~61 (
	.dataa(\u0_m0_wo0_mtree_mult1_14_add_3_o[17]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_15_sub_1_o[19]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_add0_7_o[19]~60 ),
	.combout(\u0_m0_wo0_mtree_add0_7_o[20]~61_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_add0_7_o[20]~61 .lut_mask = 16'h6969;
defparam \u0_m0_wo0_mtree_add0_7_o[20]~61 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add0_7_o[20] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[20]~61_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[20]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[20] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[20] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_7_o[19] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[19]~59_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[19]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[19] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[19] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_7_o[18] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[18]~57_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[18]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[18] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[18] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_6_o[17] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_6_o[17]~53_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_6_o[17]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_6_o[17] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_6_o[17] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_7_o[17] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[17]~55_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[17]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[17] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[17] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_6_o[16] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_6_o[16]~51_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_6_o[16]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_6_o[16] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_6_o[16] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_7_o[16] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[16]~53_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[16]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[16] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[16] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_6_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_6_o[15]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_6_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_6_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_6_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_7_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[15]~51_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_6_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_6_o[14]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_6_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_6_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_6_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_7_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[14]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_6_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_6_o[13]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_6_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_6_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_6_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_7_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[13]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_6_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_6_o[12]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_6_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_6_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_6_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_7_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[12]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_6_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_6_o[11]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_6_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_6_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_6_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_7_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[11]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_6_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_6_o[10]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_6_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_6_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_6_o[10] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_7_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_7_o[10]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_7_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_7_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_7_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[10]~41 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[10]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_3_o[9]~40 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[10]~41_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[10]~42 ));
defparam \u0_m0_wo0_mtree_add1_3_o[10]~41 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_3_o[10]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[11]~43 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[11]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_3_o[10]~42 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[11]~43_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[11]~44 ));
defparam \u0_m0_wo0_mtree_add1_3_o[11]~43 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_3_o[11]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[12]~45 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[12]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_3_o[11]~44 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[12]~45_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[12]~46 ));
defparam \u0_m0_wo0_mtree_add1_3_o[12]~45 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_3_o[12]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[13]~47 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[13]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_3_o[12]~46 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[13]~47_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[13]~48 ));
defparam \u0_m0_wo0_mtree_add1_3_o[13]~47 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_3_o[13]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[14]~49 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[14]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_3_o[13]~48 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[14]~49_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[14]~50 ));
defparam \u0_m0_wo0_mtree_add1_3_o[14]~49 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_3_o[14]~49 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[15]~51 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_3_o[14]~50 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[15]~51_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[15]~52 ));
defparam \u0_m0_wo0_mtree_add1_3_o[15]~51 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_3_o[15]~51 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[16]~53 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[16]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_3_o[15]~52 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[16]~53_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[16]~54 ));
defparam \u0_m0_wo0_mtree_add1_3_o[16]~53 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_3_o[16]~53 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[17]~55 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[17]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_3_o[16]~54 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[17]~55_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[17]~56 ));
defparam \u0_m0_wo0_mtree_add1_3_o[17]~55 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_3_o[17]~55 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[18]~57 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[18]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[18]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_3_o[17]~56 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[18]~57_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[18]~58 ));
defparam \u0_m0_wo0_mtree_add1_3_o[18]~57 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_3_o[18]~57 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[19]~59 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[18]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[19]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_3_o[18]~58 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[19]~59_combout ),
	.cout(\u0_m0_wo0_mtree_add1_3_o[19]~60 ));
defparam \u0_m0_wo0_mtree_add1_3_o[19]~59 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_3_o[19]~59 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_3_o[20]~61 (
	.dataa(\u0_m0_wo0_mtree_add0_6_o[18]~q ),
	.datab(\u0_m0_wo0_mtree_add0_7_o[20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_add1_3_o[19]~60 ),
	.combout(\u0_m0_wo0_mtree_add1_3_o[20]~61_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_add1_3_o[20]~61 .lut_mask = 16'h6969;
defparam \u0_m0_wo0_mtree_add1_3_o[20]~61 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add1_3_o[20] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[20]~61_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[20]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[20] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[20] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_3_o[19] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[19]~59_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[19]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[19] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[19] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_3_o[18] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[18]~57_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[18]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[18] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[18] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_3_o[17] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[17]~55_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[17]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[17] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[17] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_3_o[16] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[16]~53_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[16]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[16] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[16] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_2_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_2_o[15]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_2_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_2_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_2_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_3_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[15]~51_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_2_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_2_o[14]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_2_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_2_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_2_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_3_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[14]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_2_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_2_o[13]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_2_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_2_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_2_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_3_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[13]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_2_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_2_o[12]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_2_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_2_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_2_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_3_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[12]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_2_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_2_o[11]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_2_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_2_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_2_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_3_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[11]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_2_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_2_o[10]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_2_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_2_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_2_o[10] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_3_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_3_o[10]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_3_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_3_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_3_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[10]~41 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[10]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_1_o[9]~40 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[10]~41_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[10]~42 ));
defparam \u0_m0_wo0_mtree_add2_1_o[10]~41 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add2_1_o[10]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[11]~43 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[11]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_1_o[10]~42 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[11]~43_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[11]~44 ));
defparam \u0_m0_wo0_mtree_add2_1_o[11]~43 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_1_o[11]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[12]~45 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[12]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_1_o[11]~44 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[12]~45_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[12]~46 ));
defparam \u0_m0_wo0_mtree_add2_1_o[12]~45 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add2_1_o[12]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[13]~47 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[13]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_1_o[12]~46 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[13]~47_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[13]~48 ));
defparam \u0_m0_wo0_mtree_add2_1_o[13]~47 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_1_o[13]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[14]~49 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[14]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_1_o[13]~48 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[14]~49_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[14]~50 ));
defparam \u0_m0_wo0_mtree_add2_1_o[14]~49 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add2_1_o[14]~49 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[15]~51 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_1_o[14]~50 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[15]~51_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[15]~52 ));
defparam \u0_m0_wo0_mtree_add2_1_o[15]~51 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_1_o[15]~51 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[16]~53 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[17]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_1_o[15]~52 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[16]~53_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[16]~54 ));
defparam \u0_m0_wo0_mtree_add2_1_o[16]~53 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add2_1_o[16]~53 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[17]~55 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[17]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_1_o[16]~54 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[17]~55_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[17]~56 ));
defparam \u0_m0_wo0_mtree_add2_1_o[17]~55 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_1_o[17]~55 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[18]~57 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[17]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[18]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_1_o[17]~56 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[18]~57_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[18]~58 ));
defparam \u0_m0_wo0_mtree_add2_1_o[18]~57 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add2_1_o[18]~57 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[19]~59 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[17]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[19]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_1_o[18]~58 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[19]~59_combout ),
	.cout(\u0_m0_wo0_mtree_add2_1_o[19]~60 ));
defparam \u0_m0_wo0_mtree_add2_1_o[19]~59 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_1_o[19]~59 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_1_o[20]~61 (
	.dataa(\u0_m0_wo0_mtree_add1_2_o[17]~q ),
	.datab(\u0_m0_wo0_mtree_add1_3_o[20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_add2_1_o[19]~60 ),
	.combout(\u0_m0_wo0_mtree_add2_1_o[20]~61_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_add2_1_o[20]~61 .lut_mask = 16'h6969;
defparam \u0_m0_wo0_mtree_add2_1_o[20]~61 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add2_1_o[20] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[20]~61_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[20]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[20] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[20] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_1_o[19] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[19]~59_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[19]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[19] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[19] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_1_o[18] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[18]~57_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[18]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[18] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[18] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_1_o[17] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[17]~55_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[17]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[17] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[17] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_1_o[16] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[16]~53_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[16]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[16] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[16] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_1_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[15]~51_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_1_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[14]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_1_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[13]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_1_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_1_o[12]~38_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_1_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_1_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_1_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_1_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[12]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_1_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_1_o[11]~36_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_1_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_1_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_1_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_1_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[11]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_1_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_1_o[10]~34_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_1_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_1_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_1_o[10] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_1_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_1_o[10]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_1_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_1_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[10]~41 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[10]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_0_o[9]~40 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[10]~41_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[10]~42 ));
defparam \u0_m0_wo0_mtree_add3_0_o[10]~41 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add3_0_o[10]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[11]~43 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[11]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_0_o[10]~42 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[11]~43_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[11]~44 ));
defparam \u0_m0_wo0_mtree_add3_0_o[11]~43 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_0_o[11]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[12]~45 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[12]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_0_o[11]~44 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[12]~45_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[12]~46 ));
defparam \u0_m0_wo0_mtree_add3_0_o[12]~45 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add3_0_o[12]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[13]~47 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_0_o[12]~46 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[13]~47_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[13]~48 ));
defparam \u0_m0_wo0_mtree_add3_0_o[13]~47 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_0_o[13]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[14]~49 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_0_o[13]~48 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[14]~49_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[14]~50 ));
defparam \u0_m0_wo0_mtree_add3_0_o[14]~49 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add3_0_o[14]~49 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[15]~51 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_0_o[14]~50 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[15]~51_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[15]~52 ));
defparam \u0_m0_wo0_mtree_add3_0_o[15]~51 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_0_o[15]~51 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[16]~53 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_0_o[15]~52 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[16]~53_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[16]~54 ));
defparam \u0_m0_wo0_mtree_add3_0_o[16]~53 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add3_0_o[16]~53 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[17]~55 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_0_o[16]~54 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[17]~55_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[17]~56 ));
defparam \u0_m0_wo0_mtree_add3_0_o[17]~55 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_0_o[17]~55 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[18]~57 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[18]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_0_o[17]~56 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[18]~57_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[18]~58 ));
defparam \u0_m0_wo0_mtree_add3_0_o[18]~57 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add3_0_o[18]~57 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[19]~59 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[19]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_0_o[18]~58 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[19]~59_combout ),
	.cout(\u0_m0_wo0_mtree_add3_0_o[19]~60 ));
defparam \u0_m0_wo0_mtree_add3_0_o[19]~59 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_0_o[19]~59 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_0_o[20]~61 (
	.dataa(\u0_m0_wo0_mtree_add1_1_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_add2_1_o[20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_add3_0_o[19]~60 ),
	.combout(\u0_m0_wo0_mtree_add3_0_o[20]~61_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_add3_0_o[20]~61 .lut_mask = 16'h6969;
defparam \u0_m0_wo0_mtree_add3_0_o[20]~61 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add3_0_o[20] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[20]~61_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[20]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[20] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[20] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_1_o[10]~29 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][8]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_1_o[9]~28 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_1_o[10]~29_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_1_o[10]~30 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[10]~29 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[10]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_1_o[11]~31 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][9]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_1_o[10]~30 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_1_o[11]~31_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_1_o[11]~32 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[11]~31 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[11]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_1_o[12]~33 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][10]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_1_o[11]~32 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_1_o[12]~33_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_1_o[12]~34 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[12]~33 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[12]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_1_o[13]~35 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr14|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_1_o[12]~34 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_1_o[13]~35_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_1_o[13]~36 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[13]~35 .lut_mask = 16'hF0AA;
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[13]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_1_o[14]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_1_o[13]~36 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_1_o[14]~37_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[14]~37 .lut_mask = 16'hF0F0;
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[14]~37 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_16_add_1_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_1_o[14]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_1_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_1_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_1_o[13]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_1_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_1_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_1_o[12]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_1_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_1_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_1_o[11]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_1_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_1_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_1_o[10]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_1_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_3_o[10]~23 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][5]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_16_add_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_3_o[9]~22 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_3_o[10]~23_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_3_o[10]~24 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[10]~23 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[10]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_3_o[11]~25 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][6]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_16_add_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_3_o[10]~24 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_3_o[11]~25_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_3_o[11]~26 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[11]~25 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[11]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_3_o[12]~27 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][7]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_16_add_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_3_o[11]~26 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_3_o[12]~27_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_3_o[12]~28 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[12]~27 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[12]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_3_o[13]~29 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][8]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_16_add_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_3_o[12]~28 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_3_o[13]~29_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_3_o[13]~30 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[13]~29 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[13]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_3_o[14]~31 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][9]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_16_add_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_3_o[13]~30 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_3_o[14]~31_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_3_o[14]~32 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[14]~31 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[14]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_3_o[15]~33 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][10]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_16_add_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_3_o[14]~32 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_3_o[15]~33_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_3_o[15]~34 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[15]~33 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[15]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_3_o[16]~35 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_16_add_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_3_o[15]~34 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_3_o[16]~35_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_16_add_3_o[16]~36 ));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[16]~35 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[16]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_16_add_3_o[17]~37 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_16_add_1_o[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_16_add_3_o[16]~36 ),
	.combout(\u0_m0_wo0_mtree_mult1_16_add_3_o[17]~37_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[17]~37 .lut_mask = 16'h6969;
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[17]~37 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_16_add_3_o[17] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_3_o[17]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_3_o[17]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[17] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[17] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_1_o[10]~33 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][7]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_1_o[9]~32 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[10]~33_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[10]~34 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[10]~33 .lut_mask = 16'h694D;
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[10]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_1_o[11]~35 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][8]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_1_o[10]~34 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[11]~35_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[11]~36 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[11]~35 .lut_mask = 16'h962B;
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[11]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_1_o[12]~37 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][9]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_1_o[11]~36 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[12]~37_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[12]~38 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[12]~37 .lut_mask = 16'h694D;
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[12]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_1_o[13]~39 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][10]~q ),
	.datab(\u0_m0_wo0_wi0_r0_delayr13|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_1_o[12]~38 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[13]~39_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[13]~40 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[13]~39 .lut_mask = 16'h962B;
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[13]~39 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_1_o[14]~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_1_o[13]~40 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[14]~41_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[14]~42 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[14]~41 .lut_mask = 16'h0F0F;
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[14]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_1_o[15]~43 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_1_o[14]~42 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_1_o[15]~43_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[15]~43 .lut_mask = 16'hF0F0;
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[15]~43 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_1_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[15]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_1_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_1_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[14]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_1_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_1_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[13]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_1_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_1_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[12]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_1_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_1_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[11]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_1_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_1_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_1_o[10]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_1_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_3_o[10]~23 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][5]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_3_o[9]~22 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[10]~23_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[10]~24 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[10]~23 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[10]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_3_o[11]~25 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][6]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_3_o[10]~24 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[11]~25_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[11]~26 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[11]~25 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[11]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_3_o[12]~27 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][7]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_3_o[11]~26 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[12]~27_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[12]~28 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[12]~27 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[12]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_3_o[13]~29 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][8]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_3_o[12]~28 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[13]~29_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[13]~30 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[13]~29 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[13]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_3_o[14]~31 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][9]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_3_o[13]~30 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[14]~31_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[14]~32 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[14]~31 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[14]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_3_o[15]~33 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][10]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_1_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_3_o[14]~32 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[15]~33_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[15]~34 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[15]~33 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[15]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_3_o[16]~35 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_1_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_3_o[15]~34 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[16]~35_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[16]~36 ));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[16]~35 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[16]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_17_sub_3_o[17]~37 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_1_o[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_17_sub_3_o[16]~36 ),
	.combout(\u0_m0_wo0_mtree_mult1_17_sub_3_o[17]~37_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[17]~37 .lut_mask = 16'h9696;
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[17]~37 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_3_o[17] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_3_o[17]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_3_o[17]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[17] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[17] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_3_o[16] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_3_o[16]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_3_o[16]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[16] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[16] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_3_o[16] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_3_o[16]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_3_o[16]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[16] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[16] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_3_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_3_o[15]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_3_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_3_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_3_o[15]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_3_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_3_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_3_o[14]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_3_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_3_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_3_o[14]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_3_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_3_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_3_o[13]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_3_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_3_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_3_o[13]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_3_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_3_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_3_o[12]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_3_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_3_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_3_o[12]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_3_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_3_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_3_o[11]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_3_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_3_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_3_o[11]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_3_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_16_add_3_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_16_add_3_o[10]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_16_add_3_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_16_add_3_o[10] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_17_sub_3_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_17_sub_3_o[10]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_17_sub_3_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_17_sub_3_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_8_o[10]~39 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_3_o[10]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_3_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_8_o[9]~38 ),
	.combout(\u0_m0_wo0_mtree_add0_8_o[10]~39_combout ),
	.cout(\u0_m0_wo0_mtree_add0_8_o[10]~40 ));
defparam \u0_m0_wo0_mtree_add0_8_o[10]~39 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_8_o[10]~39 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_8_o[11]~41 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_3_o[11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_3_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_8_o[10]~40 ),
	.combout(\u0_m0_wo0_mtree_add0_8_o[11]~41_combout ),
	.cout(\u0_m0_wo0_mtree_add0_8_o[11]~42 ));
defparam \u0_m0_wo0_mtree_add0_8_o[11]~41 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_8_o[11]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_8_o[12]~43 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_3_o[12]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_3_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_8_o[11]~42 ),
	.combout(\u0_m0_wo0_mtree_add0_8_o[12]~43_combout ),
	.cout(\u0_m0_wo0_mtree_add0_8_o[12]~44 ));
defparam \u0_m0_wo0_mtree_add0_8_o[12]~43 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_8_o[12]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_8_o[13]~45 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_3_o[13]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_3_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_8_o[12]~44 ),
	.combout(\u0_m0_wo0_mtree_add0_8_o[13]~45_combout ),
	.cout(\u0_m0_wo0_mtree_add0_8_o[13]~46 ));
defparam \u0_m0_wo0_mtree_add0_8_o[13]~45 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_8_o[13]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_8_o[14]~47 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_3_o[14]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_3_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_8_o[13]~46 ),
	.combout(\u0_m0_wo0_mtree_add0_8_o[14]~47_combout ),
	.cout(\u0_m0_wo0_mtree_add0_8_o[14]~48 ));
defparam \u0_m0_wo0_mtree_add0_8_o[14]~47 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_8_o[14]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_8_o[15]~49 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_3_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_3_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_8_o[14]~48 ),
	.combout(\u0_m0_wo0_mtree_add0_8_o[15]~49_combout ),
	.cout(\u0_m0_wo0_mtree_add0_8_o[15]~50 ));
defparam \u0_m0_wo0_mtree_add0_8_o[15]~49 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_8_o[15]~49 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_8_o[16]~51 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_3_o[16]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_3_o[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_8_o[15]~50 ),
	.combout(\u0_m0_wo0_mtree_add0_8_o[16]~51_combout ),
	.cout(\u0_m0_wo0_mtree_add0_8_o[16]~52 ));
defparam \u0_m0_wo0_mtree_add0_8_o[16]~51 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_8_o[16]~51 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_8_o[17]~53 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_3_o[17]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_3_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_8_o[16]~52 ),
	.combout(\u0_m0_wo0_mtree_add0_8_o[17]~53_combout ),
	.cout(\u0_m0_wo0_mtree_add0_8_o[17]~54 ));
defparam \u0_m0_wo0_mtree_add0_8_o[17]~53 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_8_o[17]~53 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_8_o[18]~55 (
	.dataa(\u0_m0_wo0_mtree_mult1_16_add_3_o[17]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_17_sub_3_o[17]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_add0_8_o[17]~54 ),
	.combout(\u0_m0_wo0_mtree_add0_8_o[18]~55_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_add0_8_o[18]~55 .lut_mask = 16'h6969;
defparam \u0_m0_wo0_mtree_add0_8_o[18]~55 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add0_8_o[18] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_8_o[18]~55_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_8_o[18]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_8_o[18] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_8_o[18] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_1_o[10]~31 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][10]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_1_o[9]~30 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_1_o[10]~31_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_1_o[10]~32 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[10]~31 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[10]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_1_o[11]~33 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][10]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_1_o[10]~32 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_1_o[11]~33_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_1_o[11]~34 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[11]~33 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[11]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_1_o[12]~35 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_1_o[11]~34 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_1_o[12]~35_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_1_o[12]~36 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[12]~35 .lut_mask = 16'hF0AA;
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[12]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_1_o[13]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_1_o[12]~36 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_1_o[13]~37_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[13]~37 .lut_mask = 16'hF0F0;
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[13]~37 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_18_add_1_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_1_o[13]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_1_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_1_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_1_o[12]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_1_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_1_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_1_o[11]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_1_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_1_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_1_o[10]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_1_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_3_o[10]~27 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][7]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_3_o[9]~26 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_3_o[10]~27_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_3_o[10]~28 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[10]~27 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[10]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_3_o[11]~29 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][8]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_3_o[10]~28 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_3_o[11]~29_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_3_o[11]~30 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[11]~29 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[11]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_3_o[12]~31 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][9]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_3_o[11]~30 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_3_o[12]~31_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_3_o[12]~32 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[12]~31 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[12]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_3_o[13]~33 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][10]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_3_o[12]~32 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_3_o[13]~33_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_3_o[13]~34 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[13]~33 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[13]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_3_o[14]~35 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_3_o[13]~34 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_3_o[14]~35_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_18_add_3_o[14]~36 ));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[14]~35 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[14]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_18_add_3_o[15]~37 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_1_o[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_18_add_3_o[14]~36 ),
	.combout(\u0_m0_wo0_mtree_mult1_18_add_3_o[15]~37_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[15]~37 .lut_mask = 16'h6969;
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[15]~37 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_18_add_3_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_3_o[15]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_3_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_8_o[17] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_8_o[17]~53_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_8_o[17]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_8_o[17] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_8_o[17] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_8_o[16] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_8_o[16]~51_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_8_o[16]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_8_o[16] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_8_o[16] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_8_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_8_o[15]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_8_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_8_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_8_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_8_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_8_o[14]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_8_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_8_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_8_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_3_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_3_o[14]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_3_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_8_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_8_o[13]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_8_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_8_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_8_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_3_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_3_o[13]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_3_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_8_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_8_o[12]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_8_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_8_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_8_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_3_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_3_o[12]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_3_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_8_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_8_o[11]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_8_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_8_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_8_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_3_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_3_o[11]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_3_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_8_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_8_o[10]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_8_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_8_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_8_o[10] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_18_add_3_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_18_add_3_o[10]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_18_add_3_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_18_add_3_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[10]~40 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[10]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_4_o[9]~39 ),
	.combout(\u0_m0_wo0_mtree_add1_4_o[10]~40_combout ),
	.cout(\u0_m0_wo0_mtree_add1_4_o[10]~41 ));
defparam \u0_m0_wo0_mtree_add1_4_o[10]~40 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_4_o[10]~40 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[11]~42 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_4_o[10]~41 ),
	.combout(\u0_m0_wo0_mtree_add1_4_o[11]~42_combout ),
	.cout(\u0_m0_wo0_mtree_add1_4_o[11]~43 ));
defparam \u0_m0_wo0_mtree_add1_4_o[11]~42 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_4_o[11]~42 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[12]~44 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[12]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_4_o[11]~43 ),
	.combout(\u0_m0_wo0_mtree_add1_4_o[12]~44_combout ),
	.cout(\u0_m0_wo0_mtree_add1_4_o[12]~45 ));
defparam \u0_m0_wo0_mtree_add1_4_o[12]~44 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_4_o[12]~44 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[13]~46 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[13]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_4_o[12]~45 ),
	.combout(\u0_m0_wo0_mtree_add1_4_o[13]~46_combout ),
	.cout(\u0_m0_wo0_mtree_add1_4_o[13]~47 ));
defparam \u0_m0_wo0_mtree_add1_4_o[13]~46 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_4_o[13]~46 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[14]~48 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[14]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_4_o[13]~47 ),
	.combout(\u0_m0_wo0_mtree_add1_4_o[14]~48_combout ),
	.cout(\u0_m0_wo0_mtree_add1_4_o[14]~49 ));
defparam \u0_m0_wo0_mtree_add1_4_o[14]~48 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_4_o[14]~48 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[15]~50 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_4_o[14]~49 ),
	.combout(\u0_m0_wo0_mtree_add1_4_o[15]~50_combout ),
	.cout(\u0_m0_wo0_mtree_add1_4_o[15]~51 ));
defparam \u0_m0_wo0_mtree_add1_4_o[15]~50 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_4_o[15]~50 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[16]~52 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[16]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_4_o[15]~51 ),
	.combout(\u0_m0_wo0_mtree_add1_4_o[16]~52_combout ),
	.cout(\u0_m0_wo0_mtree_add1_4_o[16]~53 ));
defparam \u0_m0_wo0_mtree_add1_4_o[16]~52 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_4_o[16]~52 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[17]~54 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[17]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_4_o[16]~53 ),
	.combout(\u0_m0_wo0_mtree_add1_4_o[17]~54_combout ),
	.cout(\u0_m0_wo0_mtree_add1_4_o[17]~55 ));
defparam \u0_m0_wo0_mtree_add1_4_o[17]~54 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_4_o[17]~54 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[18]~56 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[18]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_4_o[17]~55 ),
	.combout(\u0_m0_wo0_mtree_add1_4_o[18]~56_combout ),
	.cout(\u0_m0_wo0_mtree_add1_4_o[18]~57 ));
defparam \u0_m0_wo0_mtree_add1_4_o[18]~56 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_4_o[18]~56 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_4_o[20]~58 (
	.dataa(\u0_m0_wo0_mtree_add0_8_o[18]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_18_add_3_o[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_add1_4_o[18]~57 ),
	.combout(\u0_m0_wo0_mtree_add1_4_o[20]~58_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_add1_4_o[20]~58 .lut_mask = 16'h9696;
defparam \u0_m0_wo0_mtree_add1_4_o[20]~58 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add1_4_o[20] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[20]~58_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[20]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[20] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[20] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_0_o[10]~30 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_0_o[9]~29 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[10]~30_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[10]~31 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[10]~30 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[10]~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_0_o[11]~32 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_0_o[10]~31 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[11]~32_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[11]~33 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[11]~32 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[11]~32 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_0_o[12]~34 (
	.dataa(\u0_m0_wo0_wi0_r0_delayr10|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_0_o[11]~33 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_0_o[12]~34_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[12]~34 .lut_mask = 16'hA5A5;
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[12]~34 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_0_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_0_o[12]~34_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_0_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_0_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_0_o[11]~32_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_0_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_0_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_0_o[10]~30_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_0_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_0_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_2_o[10]~29 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][8]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_20_sub_0_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_2_o[9]~28 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[10]~29_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[10]~30 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[10]~29 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[10]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_2_o[11]~31 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][9]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_20_sub_0_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_2_o[10]~30 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[11]~31_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[11]~32 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[11]~31 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[11]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_2_o[12]~33 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][10]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_20_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_2_o[11]~32 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[12]~33_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[12]~34 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[12]~33 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[12]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_2_o[13]~35 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_20_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_2_o[12]~34 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[13]~35_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[13]~36 ));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[13]~35 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[13]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_20_sub_2_o[14]~37 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_20_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_20_sub_2_o[13]~36 ),
	.combout(\u0_m0_wo0_mtree_mult1_20_sub_2_o[14]~37_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[14]~37 .lut_mask = 16'h9696;
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[14]~37 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_2_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_2_o[14]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_2_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[14] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_21_add_1_o[9]~29 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][8]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_21_add_1_o[8]~28 ),
	.combout(\u0_m0_wo0_mtree_mult1_21_add_1_o[9]~29_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_21_add_1_o[9]~30 ));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[9]~29 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[9]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_21_add_1_o[10]~31 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][10]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_21_add_1_o[9]~30 ),
	.combout(\u0_m0_wo0_mtree_mult1_21_add_1_o[10]~31_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_21_add_1_o[10]~32 ));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[10]~31 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[10]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_21_add_1_o[11]~33 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][10]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_21_add_1_o[10]~32 ),
	.combout(\u0_m0_wo0_mtree_mult1_21_add_1_o[11]~33_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_21_add_1_o[11]~34 ));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[11]~33 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[11]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_21_add_1_o[12]~35 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_21_add_1_o[11]~34 ),
	.combout(\u0_m0_wo0_mtree_mult1_21_add_1_o[12]~35_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_21_add_1_o[12]~36 ));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[12]~35 .lut_mask = 16'hF0AA;
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[12]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_21_add_1_o[13]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_21_add_1_o[12]~36 ),
	.combout(\u0_m0_wo0_mtree_mult1_21_add_1_o[13]~37_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[13]~37 .lut_mask = 16'hF0F0;
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[13]~37 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_21_add_1_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_21_add_1_o[13]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_21_add_1_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_2_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_2_o[13]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_2_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_21_add_1_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_21_add_1_o[12]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_21_add_1_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_2_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_2_o[12]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_2_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_21_add_1_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_21_add_1_o[11]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_21_add_1_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_2_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_2_o[11]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_2_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_21_add_1_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_21_add_1_o[10]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_21_add_1_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[10] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_20_sub_2_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_20_sub_2_o[10]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_20_sub_2_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_20_sub_2_o[10] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_21_add_1_o[9] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_21_add_1_o[9]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_21_add_1_o[9]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[9] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_21_add_1_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_10_o[10]~33 (
	.dataa(\u0_m0_wo0_mtree_mult1_20_sub_2_o[10]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_21_add_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_10_o[9]~32 ),
	.combout(\u0_m0_wo0_mtree_add0_10_o[10]~33_combout ),
	.cout(\u0_m0_wo0_mtree_add0_10_o[10]~34 ));
defparam \u0_m0_wo0_mtree_add0_10_o[10]~33 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_10_o[10]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_10_o[11]~35 (
	.dataa(\u0_m0_wo0_mtree_mult1_20_sub_2_o[11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_21_add_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_10_o[10]~34 ),
	.combout(\u0_m0_wo0_mtree_add0_10_o[11]~35_combout ),
	.cout(\u0_m0_wo0_mtree_add0_10_o[11]~36 ));
defparam \u0_m0_wo0_mtree_add0_10_o[11]~35 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_10_o[11]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_10_o[12]~37 (
	.dataa(\u0_m0_wo0_mtree_mult1_20_sub_2_o[12]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_21_add_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_10_o[11]~36 ),
	.combout(\u0_m0_wo0_mtree_add0_10_o[12]~37_combout ),
	.cout(\u0_m0_wo0_mtree_add0_10_o[12]~38 ));
defparam \u0_m0_wo0_mtree_add0_10_o[12]~37 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_10_o[12]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_10_o[13]~39 (
	.dataa(\u0_m0_wo0_mtree_mult1_20_sub_2_o[13]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_21_add_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_10_o[12]~38 ),
	.combout(\u0_m0_wo0_mtree_add0_10_o[13]~39_combout ),
	.cout(\u0_m0_wo0_mtree_add0_10_o[13]~40 ));
defparam \u0_m0_wo0_mtree_add0_10_o[13]~39 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_10_o[13]~39 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_10_o[14]~41 (
	.dataa(\u0_m0_wo0_mtree_mult1_20_sub_2_o[14]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_21_add_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_10_o[13]~40 ),
	.combout(\u0_m0_wo0_mtree_add0_10_o[14]~41_combout ),
	.cout(\u0_m0_wo0_mtree_add0_10_o[14]~42 ));
defparam \u0_m0_wo0_mtree_add0_10_o[14]~41 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_10_o[14]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_10_o[15]~43 (
	.dataa(\u0_m0_wo0_mtree_mult1_20_sub_2_o[14]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_21_add_1_o[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_add0_10_o[14]~42 ),
	.combout(\u0_m0_wo0_mtree_add0_10_o[15]~43_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_add0_10_o[15]~43 .lut_mask = 16'h6969;
defparam \u0_m0_wo0_mtree_add0_10_o[15]~43 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add0_10_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_10_o[15]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_10_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_10_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_10_o[15] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_22_sub_1_o[10]~29 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][8]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_22_sub_1_o[9]~28 ),
	.combout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[10]~29_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[10]~30 ));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[10]~29 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[10]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_22_sub_1_o[11]~31 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][9]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_22_sub_1_o[10]~30 ),
	.combout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[11]~31_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[11]~32 ));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[11]~31 .lut_mask = 16'h692B;
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[11]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_22_sub_1_o[12]~33 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][10]~q ),
	.datab(\d_u0_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_22_sub_1_o[11]~32 ),
	.combout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[12]~33_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[12]~34 ));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[12]~33 .lut_mask = 16'h964D;
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[12]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_22_sub_1_o[13]~35 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_22_sub_1_o[12]~34 ),
	.combout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[13]~35_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[13]~36 ));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[13]~35 .lut_mask = 16'h0F0F;
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[13]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_22_sub_1_o[14]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_22_sub_1_o[13]~36 ),
	.combout(\u0_m0_wo0_mtree_mult1_22_sub_1_o[14]~37_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[14]~37 .lut_mask = 16'hF0F0;
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[14]~37 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_22_sub_1_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_22_sub_1_o[14]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_22_sub_1_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_10_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_10_o[14]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_10_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_10_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_10_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_10_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_10_o[13]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_10_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_10_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_10_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_22_sub_1_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_22_sub_1_o[13]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_22_sub_1_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_10_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_10_o[12]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_10_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_10_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_10_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_22_sub_1_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_22_sub_1_o[12]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_22_sub_1_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_10_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_10_o[11]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_10_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_10_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_10_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_22_sub_1_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_22_sub_1_o[11]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_22_sub_1_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_10_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_10_o[10]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_10_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_10_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_10_o[10] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_22_sub_1_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_22_sub_1_o[10]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_22_sub_1_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_22_sub_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_5_o[10]~37 (
	.dataa(\u0_m0_wo0_mtree_add0_10_o[10]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_22_sub_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_5_o[9]~36 ),
	.combout(\u0_m0_wo0_mtree_add1_5_o[10]~37_combout ),
	.cout(\u0_m0_wo0_mtree_add1_5_o[10]~38 ));
defparam \u0_m0_wo0_mtree_add1_5_o[10]~37 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_5_o[10]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_5_o[11]~39 (
	.dataa(\u0_m0_wo0_mtree_add0_10_o[11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_22_sub_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_5_o[10]~38 ),
	.combout(\u0_m0_wo0_mtree_add1_5_o[11]~39_combout ),
	.cout(\u0_m0_wo0_mtree_add1_5_o[11]~40 ));
defparam \u0_m0_wo0_mtree_add1_5_o[11]~39 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_5_o[11]~39 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_5_o[12]~41 (
	.dataa(\u0_m0_wo0_mtree_add0_10_o[12]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_22_sub_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_5_o[11]~40 ),
	.combout(\u0_m0_wo0_mtree_add1_5_o[12]~41_combout ),
	.cout(\u0_m0_wo0_mtree_add1_5_o[12]~42 ));
defparam \u0_m0_wo0_mtree_add1_5_o[12]~41 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_5_o[12]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_5_o[13]~43 (
	.dataa(\u0_m0_wo0_mtree_add0_10_o[13]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_22_sub_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_5_o[12]~42 ),
	.combout(\u0_m0_wo0_mtree_add1_5_o[13]~43_combout ),
	.cout(\u0_m0_wo0_mtree_add1_5_o[13]~44 ));
defparam \u0_m0_wo0_mtree_add1_5_o[13]~43 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_5_o[13]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_5_o[14]~45 (
	.dataa(\u0_m0_wo0_mtree_add0_10_o[14]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_22_sub_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_5_o[13]~44 ),
	.combout(\u0_m0_wo0_mtree_add1_5_o[14]~45_combout ),
	.cout(\u0_m0_wo0_mtree_add1_5_o[14]~46 ));
defparam \u0_m0_wo0_mtree_add1_5_o[14]~45 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add1_5_o[14]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_5_o[15]~47 (
	.dataa(\u0_m0_wo0_mtree_add0_10_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_22_sub_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add1_5_o[14]~46 ),
	.combout(\u0_m0_wo0_mtree_add1_5_o[15]~47_combout ),
	.cout(\u0_m0_wo0_mtree_add1_5_o[15]~48 ));
defparam \u0_m0_wo0_mtree_add1_5_o[15]~47 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add1_5_o[15]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add1_5_o[17]~49 (
	.dataa(\u0_m0_wo0_mtree_add0_10_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_22_sub_1_o[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_add1_5_o[15]~48 ),
	.combout(\u0_m0_wo0_mtree_add1_5_o[17]~49_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_add1_5_o[17]~49 .lut_mask = 16'h6969;
defparam \u0_m0_wo0_mtree_add1_5_o[17]~49 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add1_5_o[17] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_5_o[17]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_5_o[17]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_5_o[17] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_5_o[17] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_4_o[18] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[18]~56_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[18]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[18] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[18] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_4_o[17] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[17]~54_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[17]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[17] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[17] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_4_o[16] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[16]~52_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[16]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[16] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[16] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_4_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[15]~50_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_5_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_5_o[15]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_5_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_5_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_5_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_4_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[14]~48_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_5_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_5_o[14]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_5_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_5_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_5_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_4_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[13]~46_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_5_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_5_o[13]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_5_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_5_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_5_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_4_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[12]~44_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_5_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_5_o[12]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_5_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_5_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_5_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_4_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[11]~42_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_5_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_5_o[11]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_5_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_5_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_5_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_4_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_4_o[10]~40_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_4_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_4_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_4_o[10] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add1_5_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add1_5_o[10]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add1_5_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add1_5_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add1_5_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[10]~41 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[10]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_2_o[9]~40 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[10]~41_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[10]~42 ));
defparam \u0_m0_wo0_mtree_add2_2_o[10]~41 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add2_2_o[10]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[11]~43 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[11]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_2_o[10]~42 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[11]~43_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[11]~44 ));
defparam \u0_m0_wo0_mtree_add2_2_o[11]~43 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_2_o[11]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[12]~45 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[12]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_2_o[11]~44 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[12]~45_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[12]~46 ));
defparam \u0_m0_wo0_mtree_add2_2_o[12]~45 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add2_2_o[12]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[13]~47 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[13]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_2_o[12]~46 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[13]~47_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[13]~48 ));
defparam \u0_m0_wo0_mtree_add2_2_o[13]~47 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_2_o[13]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[14]~49 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[14]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_2_o[13]~48 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[14]~49_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[14]~50 ));
defparam \u0_m0_wo0_mtree_add2_2_o[14]~49 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add2_2_o[14]~49 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[15]~51 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_2_o[14]~50 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[15]~51_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[15]~52 ));
defparam \u0_m0_wo0_mtree_add2_2_o[15]~51 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_2_o[15]~51 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[16]~53 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[16]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_2_o[15]~52 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[16]~53_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[16]~54 ));
defparam \u0_m0_wo0_mtree_add2_2_o[16]~53 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add2_2_o[16]~53 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[17]~55 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[17]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_2_o[16]~54 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[17]~55_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[17]~56 ));
defparam \u0_m0_wo0_mtree_add2_2_o[17]~55 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_2_o[17]~55 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[18]~57 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[18]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_2_o[17]~56 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[18]~57_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[18]~58 ));
defparam \u0_m0_wo0_mtree_add2_2_o[18]~57 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add2_2_o[18]~57 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[19]~59 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[20]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add2_2_o[18]~58 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[19]~59_combout ),
	.cout(\u0_m0_wo0_mtree_add2_2_o[19]~60 ));
defparam \u0_m0_wo0_mtree_add2_2_o[19]~59 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add2_2_o[19]~59 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add2_2_o[20]~61 (
	.dataa(\u0_m0_wo0_mtree_add1_4_o[20]~q ),
	.datab(\u0_m0_wo0_mtree_add1_5_o[17]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_add2_2_o[19]~60 ),
	.combout(\u0_m0_wo0_mtree_add2_2_o[20]~61_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_add2_2_o[20]~61 .lut_mask = 16'h6969;
defparam \u0_m0_wo0_mtree_add2_2_o[20]~61 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add2_2_o[20] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[20]~61_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[20]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[20] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[20] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_25_sub_0_o[10]~30 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_25_sub_0_o[9]~29 ),
	.combout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[10]~30_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[10]~31 ));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[10]~30 .lut_mask = 16'hA5AF;
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[10]~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_25_sub_0_o[11]~32 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_mult1_25_sub_0_o[10]~31 ),
	.combout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[11]~32_combout ),
	.cout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[11]~33 ));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[11]~32 .lut_mask = 16'h5A05;
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[11]~32 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_mult1_25_sub_0_o[12]~34 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_mult1_25_sub_0_o[11]~33 ),
	.combout(\u0_m0_wo0_mtree_mult1_25_sub_0_o[12]~34_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[12]~34 .lut_mask = 16'hA5A5;
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[12]~34 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_mult1_25_sub_0_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_25_sub_0_o[12]~34_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_25_sub_0_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_25_sub_0_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_25_sub_0_o[11]~32_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_25_sub_0_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_mult1_25_sub_0_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_mult1_25_sub_0_o[10]~30_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_mult1_25_sub_0_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_mult1_25_sub_0_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_12_o[10]~34 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][10]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_25_sub_0_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_12_o[9]~33 ),
	.combout(\u0_m0_wo0_mtree_add0_12_o[10]~34_combout ),
	.cout(\u0_m0_wo0_mtree_add0_12_o[10]~35 ));
defparam \u0_m0_wo0_mtree_add0_12_o[10]~34 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_12_o[10]~34 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_12_o[11]~36 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_25_sub_0_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_12_o[10]~35 ),
	.combout(\u0_m0_wo0_mtree_add0_12_o[11]~36_combout ),
	.cout(\u0_m0_wo0_mtree_add0_12_o[11]~37 ));
defparam \u0_m0_wo0_mtree_add0_12_o[11]~36 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add0_12_o[11]~36 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_12_o[12]~38 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_25_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add0_12_o[11]~37 ),
	.combout(\u0_m0_wo0_mtree_add0_12_o[12]~38_combout ),
	.cout(\u0_m0_wo0_mtree_add0_12_o[12]~39 ));
defparam \u0_m0_wo0_mtree_add0_12_o[12]~38 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add0_12_o[12]~38 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add0_12_o[13]~40 (
	.dataa(\d_u0_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][11]~q ),
	.datab(\u0_m0_wo0_mtree_mult1_25_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_add0_12_o[12]~39 ),
	.combout(\u0_m0_wo0_mtree_add0_12_o[13]~40_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_add0_12_o[13]~40 .lut_mask = 16'h9696;
defparam \u0_m0_wo0_mtree_add0_12_o[13]~40 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add0_12_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_12_o[13]~40_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_12_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_12_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_12_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_2_o[19] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[19]~59_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[19]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[19] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[19] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_2_o[18] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[18]~57_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[18]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[18] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[18] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_2_o[17] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[17]~55_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[17]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[17] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[17] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_2_o[16] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[16]~53_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[16]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[16] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[16] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_2_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[15]~51_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_2_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[14]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_2_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[13]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_2_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[12]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_12_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_12_o[12]~38_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_12_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_12_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_12_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_2_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[11]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_12_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_12_o[11]~36_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_12_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_12_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_12_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add2_2_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add2_2_o[10]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add2_2_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add2_2_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add2_2_o[10] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add0_12_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add0_12_o[10]~34_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add0_12_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add0_12_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add0_12_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[10]~41 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[10]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_1_o[9]~40 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[10]~41_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[10]~42 ));
defparam \u0_m0_wo0_mtree_add3_1_o[10]~41 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add3_1_o[10]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[11]~43 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[11]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_1_o[10]~42 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[11]~43_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[11]~44 ));
defparam \u0_m0_wo0_mtree_add3_1_o[11]~43 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_1_o[11]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[12]~45 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[12]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_1_o[11]~44 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[12]~45_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[12]~46 ));
defparam \u0_m0_wo0_mtree_add3_1_o[12]~45 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add3_1_o[12]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[13]~47 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[13]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_1_o[12]~46 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[13]~47_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[13]~48 ));
defparam \u0_m0_wo0_mtree_add3_1_o[13]~47 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_1_o[13]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[14]~49 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[14]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_1_o[13]~48 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[14]~49_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[14]~50 ));
defparam \u0_m0_wo0_mtree_add3_1_o[14]~49 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add3_1_o[14]~49 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[15]~51 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_1_o[14]~50 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[15]~51_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[15]~52 ));
defparam \u0_m0_wo0_mtree_add3_1_o[15]~51 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_1_o[15]~51 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[16]~53 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[16]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_1_o[15]~52 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[16]~53_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[16]~54 ));
defparam \u0_m0_wo0_mtree_add3_1_o[16]~53 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add3_1_o[16]~53 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[17]~55 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[17]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_1_o[16]~54 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[17]~55_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[17]~56 ));
defparam \u0_m0_wo0_mtree_add3_1_o[17]~55 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_1_o[17]~55 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[18]~57 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[18]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_1_o[17]~56 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[18]~57_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[18]~58 ));
defparam \u0_m0_wo0_mtree_add3_1_o[18]~57 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add3_1_o[18]~57 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[19]~59 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[19]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add3_1_o[18]~58 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[19]~59_combout ),
	.cout(\u0_m0_wo0_mtree_add3_1_o[19]~60 ));
defparam \u0_m0_wo0_mtree_add3_1_o[19]~59 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add3_1_o[19]~59 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add3_1_o[20]~61 (
	.dataa(\u0_m0_wo0_mtree_add2_2_o[20]~q ),
	.datab(\u0_m0_wo0_mtree_add0_12_o[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_add3_1_o[19]~60 ),
	.combout(\u0_m0_wo0_mtree_add3_1_o[20]~61_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_add3_1_o[20]~61 .lut_mask = 16'h6969;
defparam \u0_m0_wo0_mtree_add3_1_o[20]~61 .sum_lutc_input = "cin";

dffeas \u0_m0_wo0_mtree_add3_1_o[20] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[20]~61_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[20]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[20] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[20] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_0_o[19] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[19]~59_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[19]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[19] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[19] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_1_o[19] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[19]~59_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[19]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[19] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[19] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_0_o[18] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[18]~57_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[18]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[18] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[18] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_1_o[18] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[18]~57_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[18]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[18] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[18] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_0_o[17] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[17]~55_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[17]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[17] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[17] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_1_o[17] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[17]~55_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[17]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[17] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[17] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_0_o[16] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[16]~53_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[16]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[16] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[16] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_1_o[16] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[16]~53_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[16]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[16] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[16] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_0_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[15]~51_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_1_o[15] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[15]~51_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[15]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[15] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[15] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_0_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[14]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_1_o[14] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[14]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[14]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[14] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[14] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_0_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[13]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_1_o[13] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[13]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[13]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[13] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[13] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_0_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[12]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_1_o[12] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[12]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[12]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[12] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[12] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_0_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[11]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_1_o[11] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[11]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[11]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[11] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[11] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_0_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_0_o[10]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_0_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_0_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_0_o[10] .power_up = "low";

dffeas \u0_m0_wo0_mtree_add3_1_o[10] (
	.clk(clk),
	.d(\u0_m0_wo0_mtree_add3_1_o[10]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u0_m0_wo0_mtree_add3_1_o[10]~q ),
	.prn(vcc));
defparam \u0_m0_wo0_mtree_add3_1_o[10] .is_wysiwyg = "true";
defparam \u0_m0_wo0_mtree_add3_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[10]~32 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[10]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add4_0_o[9]~31 ),
	.combout(\u0_m0_wo0_mtree_add4_0_o[10]~32_combout ),
	.cout(\u0_m0_wo0_mtree_add4_0_o[10]~33 ));
defparam \u0_m0_wo0_mtree_add4_0_o[10]~32 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add4_0_o[10]~32 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[11]~34 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[11]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add4_0_o[10]~33 ),
	.combout(\u0_m0_wo0_mtree_add4_0_o[11]~34_combout ),
	.cout(\u0_m0_wo0_mtree_add4_0_o[11]~35 ));
defparam \u0_m0_wo0_mtree_add4_0_o[11]~34 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add4_0_o[11]~34 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[12]~36 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[12]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add4_0_o[11]~35 ),
	.combout(\u0_m0_wo0_mtree_add4_0_o[12]~36_combout ),
	.cout(\u0_m0_wo0_mtree_add4_0_o[12]~37 ));
defparam \u0_m0_wo0_mtree_add4_0_o[12]~36 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add4_0_o[12]~36 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[13]~38 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[13]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add4_0_o[12]~37 ),
	.combout(\u0_m0_wo0_mtree_add4_0_o[13]~38_combout ),
	.cout(\u0_m0_wo0_mtree_add4_0_o[13]~39 ));
defparam \u0_m0_wo0_mtree_add4_0_o[13]~38 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add4_0_o[13]~38 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[14]~40 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[14]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add4_0_o[13]~39 ),
	.combout(\u0_m0_wo0_mtree_add4_0_o[14]~40_combout ),
	.cout(\u0_m0_wo0_mtree_add4_0_o[14]~41 ));
defparam \u0_m0_wo0_mtree_add4_0_o[14]~40 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add4_0_o[14]~40 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[15]~42 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[15]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add4_0_o[14]~41 ),
	.combout(\u0_m0_wo0_mtree_add4_0_o[15]~42_combout ),
	.cout(\u0_m0_wo0_mtree_add4_0_o[15]~43 ));
defparam \u0_m0_wo0_mtree_add4_0_o[15]~42 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add4_0_o[15]~42 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[16]~44 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[16]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add4_0_o[15]~43 ),
	.combout(\u0_m0_wo0_mtree_add4_0_o[16]~44_combout ),
	.cout(\u0_m0_wo0_mtree_add4_0_o[16]~45 ));
defparam \u0_m0_wo0_mtree_add4_0_o[16]~44 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add4_0_o[16]~44 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[17]~46 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[17]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add4_0_o[16]~45 ),
	.combout(\u0_m0_wo0_mtree_add4_0_o[17]~46_combout ),
	.cout(\u0_m0_wo0_mtree_add4_0_o[17]~47 ));
defparam \u0_m0_wo0_mtree_add4_0_o[17]~46 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add4_0_o[17]~46 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[18]~48 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[18]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[18]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add4_0_o[17]~47 ),
	.combout(\u0_m0_wo0_mtree_add4_0_o[18]~48_combout ),
	.cout(\u0_m0_wo0_mtree_add4_0_o[18]~49 ));
defparam \u0_m0_wo0_mtree_add4_0_o[18]~48 .lut_mask = 16'h698E;
defparam \u0_m0_wo0_mtree_add4_0_o[18]~48 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[19]~50 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[19]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[19]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u0_m0_wo0_mtree_add4_0_o[18]~49 ),
	.combout(\u0_m0_wo0_mtree_add4_0_o[19]~50_combout ),
	.cout(\u0_m0_wo0_mtree_add4_0_o[19]~51 ));
defparam \u0_m0_wo0_mtree_add4_0_o[19]~50 .lut_mask = 16'h9617;
defparam \u0_m0_wo0_mtree_add4_0_o[19]~50 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u0_m0_wo0_mtree_add4_0_o[20]~52 (
	.dataa(\u0_m0_wo0_mtree_add3_0_o[20]~q ),
	.datab(\u0_m0_wo0_mtree_add3_1_o[20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u0_m0_wo0_mtree_add4_0_o[19]~51 ),
	.combout(\u0_m0_wo0_mtree_add4_0_o[20]~52_combout ),
	.cout());
defparam \u0_m0_wo0_mtree_add4_0_o[20]~52 .lut_mask = 16'h6969;
defparam \u0_m0_wo0_mtree_add4_0_o[20]~52 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_5_sub_0_o[10]~30 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_5_sub_0_o[9]~29 ),
	.combout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[10]~30_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[10]~31 ));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[10]~30 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[10]~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_5_sub_0_o[11]~32 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_5_sub_0_o[10]~31 ),
	.combout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[11]~32_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[11]~33 ));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[11]~32 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[11]~32 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_5_sub_0_o[12]~34 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr25|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_5_sub_0_o[11]~33 ),
	.combout(\u1_m0_wo0_mtree_mult1_5_sub_0_o[12]~34_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[12]~34 .lut_mask = 16'hA5A5;
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[12]~34 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_5_sub_0_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_5_sub_0_o[12]~34_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_5_sub_0_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_5_sub_0_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_5_sub_0_o[11]~32_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_5_sub_0_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_5_sub_0_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_5_sub_0_o[10]~30_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_5_sub_0_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_5_sub_0_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_1_o[10]~34 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][10]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_5_sub_0_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_1_o[9]~33 ),
	.combout(\u1_m0_wo0_mtree_add1_1_o[10]~34_combout ),
	.cout(\u1_m0_wo0_mtree_add1_1_o[10]~35 ));
defparam \u1_m0_wo0_mtree_add1_1_o[10]~34 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_1_o[10]~34 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_1_o[11]~36 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_5_sub_0_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_1_o[10]~35 ),
	.combout(\u1_m0_wo0_mtree_add1_1_o[11]~36_combout ),
	.cout(\u1_m0_wo0_mtree_add1_1_o[11]~37 ));
defparam \u1_m0_wo0_mtree_add1_1_o[11]~36 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_1_o[11]~36 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_1_o[12]~38 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_5_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_1_o[11]~37 ),
	.combout(\u1_m0_wo0_mtree_add1_1_o[12]~38_combout ),
	.cout(\u1_m0_wo0_mtree_add1_1_o[12]~39 ));
defparam \u1_m0_wo0_mtree_add1_1_o[12]~38 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_1_o[12]~38 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_1_o[15]~40 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr24_q_14|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_5_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_add1_1_o[12]~39 ),
	.combout(\u1_m0_wo0_mtree_add1_1_o[15]~40_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_add1_1_o[15]~40 .lut_mask = 16'h9696;
defparam \u1_m0_wo0_mtree_add1_1_o[15]~40 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add1_1_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_1_o[15]~40_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_1_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_1_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_1_o[15] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_8_sub_1_o[10]~29 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][8]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_8_sub_1_o[9]~28 ),
	.combout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[10]~29_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[10]~30 ));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[10]~29 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[10]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_8_sub_1_o[11]~31 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][9]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_8_sub_1_o[10]~30 ),
	.combout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[11]~31_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[11]~32 ));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[11]~31 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[11]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_8_sub_1_o[12]~33 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][10]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr22|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_8_sub_1_o[11]~32 ),
	.combout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[12]~33_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[12]~34 ));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[12]~33 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[12]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_8_sub_1_o[13]~35 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_8_sub_1_o[12]~34 ),
	.combout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[13]~35_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[13]~36 ));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[13]~35 .lut_mask = 16'h0F0F;
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[13]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_8_sub_1_o[14]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_8_sub_1_o[13]~36 ),
	.combout(\u1_m0_wo0_mtree_mult1_8_sub_1_o[14]~37_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[14]~37 .lut_mask = 16'hF0F0;
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[14]~37 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_8_sub_1_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_8_sub_1_o[14]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_8_sub_1_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[14] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_9_add_1_o[9]~29 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][8]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_9_add_1_o[8]~28 ),
	.combout(\u1_m0_wo0_mtree_mult1_9_add_1_o[9]~29_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_9_add_1_o[9]~30 ));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[9]~29 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[9]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_9_add_1_o[10]~31 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][10]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_9_add_1_o[9]~30 ),
	.combout(\u1_m0_wo0_mtree_mult1_9_add_1_o[10]~31_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_9_add_1_o[10]~32 ));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[10]~31 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[10]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_9_add_1_o[11]~33 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][10]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_9_add_1_o[10]~32 ),
	.combout(\u1_m0_wo0_mtree_mult1_9_add_1_o[11]~33_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_9_add_1_o[11]~34 ));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[11]~33 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[11]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_9_add_1_o[12]~35 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr21|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_9_add_1_o[11]~34 ),
	.combout(\u1_m0_wo0_mtree_mult1_9_add_1_o[12]~35_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_9_add_1_o[12]~36 ));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[12]~35 .lut_mask = 16'hF0AA;
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[12]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_9_add_1_o[13]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_9_add_1_o[12]~36 ),
	.combout(\u1_m0_wo0_mtree_mult1_9_add_1_o[13]~37_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[13]~37 .lut_mask = 16'hF0F0;
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[13]~37 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_9_add_1_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_9_add_1_o[13]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_9_add_1_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_8_sub_1_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_8_sub_1_o[13]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_8_sub_1_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_9_add_1_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_9_add_1_o[12]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_9_add_1_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_8_sub_1_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_8_sub_1_o[12]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_8_sub_1_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_9_add_1_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_9_add_1_o[11]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_9_add_1_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_8_sub_1_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_8_sub_1_o[11]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_8_sub_1_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_9_add_1_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_9_add_1_o[10]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_9_add_1_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[10] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_8_sub_1_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_8_sub_1_o[10]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_8_sub_1_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_8_sub_1_o[10] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_9_add_1_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_9_add_1_o[9]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_9_add_1_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_9_add_1_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_4_o[10]~33 (
	.dataa(\u1_m0_wo0_mtree_mult1_8_sub_1_o[10]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_9_add_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_4_o[9]~32 ),
	.combout(\u1_m0_wo0_mtree_add0_4_o[10]~33_combout ),
	.cout(\u1_m0_wo0_mtree_add0_4_o[10]~34 ));
defparam \u1_m0_wo0_mtree_add0_4_o[10]~33 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_4_o[10]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_4_o[11]~35 (
	.dataa(\u1_m0_wo0_mtree_mult1_8_sub_1_o[11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_9_add_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_4_o[10]~34 ),
	.combout(\u1_m0_wo0_mtree_add0_4_o[11]~35_combout ),
	.cout(\u1_m0_wo0_mtree_add0_4_o[11]~36 ));
defparam \u1_m0_wo0_mtree_add0_4_o[11]~35 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_4_o[11]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_4_o[12]~37 (
	.dataa(\u1_m0_wo0_mtree_mult1_8_sub_1_o[12]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_9_add_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_4_o[11]~36 ),
	.combout(\u1_m0_wo0_mtree_add0_4_o[12]~37_combout ),
	.cout(\u1_m0_wo0_mtree_add0_4_o[12]~38 ));
defparam \u1_m0_wo0_mtree_add0_4_o[12]~37 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_4_o[12]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_4_o[13]~39 (
	.dataa(\u1_m0_wo0_mtree_mult1_8_sub_1_o[13]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_9_add_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_4_o[12]~38 ),
	.combout(\u1_m0_wo0_mtree_add0_4_o[13]~39_combout ),
	.cout(\u1_m0_wo0_mtree_add0_4_o[13]~40 ));
defparam \u1_m0_wo0_mtree_add0_4_o[13]~39 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_4_o[13]~39 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_4_o[14]~41 (
	.dataa(\u1_m0_wo0_mtree_mult1_8_sub_1_o[14]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_9_add_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_4_o[13]~40 ),
	.combout(\u1_m0_wo0_mtree_add0_4_o[14]~41_combout ),
	.cout(\u1_m0_wo0_mtree_add0_4_o[14]~42 ));
defparam \u1_m0_wo0_mtree_add0_4_o[14]~41 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_4_o[14]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_4_o[15]~43 (
	.dataa(\u1_m0_wo0_mtree_mult1_8_sub_1_o[14]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_9_add_1_o[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_add0_4_o[14]~42 ),
	.combout(\u1_m0_wo0_mtree_add0_4_o[15]~43_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_add0_4_o[15]~43 .lut_mask = 16'h6969;
defparam \u1_m0_wo0_mtree_add0_4_o[15]~43 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add0_4_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_4_o[15]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_4_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_4_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_4_o[15] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_0_o[10]~30 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_0_o[9]~29 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[10]~30_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[10]~31 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[10]~30 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[10]~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_0_o[11]~32 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_0_o[10]~31 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[11]~32_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[11]~33 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[11]~32 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[11]~32 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_0_o[12]~34 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr20|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_0_o[11]~33 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_0_o[12]~34_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[12]~34 .lut_mask = 16'hA5A5;
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[12]~34 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_0_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_0_o[12]~34_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_0_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_0_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_0_o[11]~32_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_0_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_0_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_0_o[10]~30_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_0_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_0_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_2_o[10]~29 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][8]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_0_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_2_o[9]~28 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[10]~29_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[10]~30 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[10]~29 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[10]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_2_o[11]~31 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][9]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_0_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_2_o[10]~30 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[11]~31_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[11]~32 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[11]~31 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[11]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_2_o[12]~33 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][10]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_2_o[11]~32 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[12]~33_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[12]~34 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[12]~33 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[12]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_2_o[13]~35 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_2_o[12]~34 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[13]~35_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[13]~36 ));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[13]~35 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[13]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_10_sub_2_o[14]~37 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr20_q_12|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_10_sub_2_o[13]~36 ),
	.combout(\u1_m0_wo0_mtree_mult1_10_sub_2_o[14]~37_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[14]~37 .lut_mask = 16'h9696;
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[14]~37 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_2_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_2_o[14]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_2_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_4_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_4_o[14]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_4_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_4_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_4_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_4_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_4_o[13]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_4_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_4_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_4_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_2_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_2_o[13]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_2_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_4_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_4_o[12]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_4_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_4_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_4_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_2_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_2_o[12]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_2_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_4_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_4_o[11]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_4_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_4_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_4_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_2_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_2_o[11]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_2_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_4_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_4_o[10]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_4_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_4_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_4_o[10] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_10_sub_2_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_10_sub_2_o[10]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_10_sub_2_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_10_sub_2_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_2_o[10]~37 (
	.dataa(\u1_m0_wo0_mtree_add0_4_o[10]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_2_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_2_o[9]~36 ),
	.combout(\u1_m0_wo0_mtree_add1_2_o[10]~37_combout ),
	.cout(\u1_m0_wo0_mtree_add1_2_o[10]~38 ));
defparam \u1_m0_wo0_mtree_add1_2_o[10]~37 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_2_o[10]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_2_o[11]~39 (
	.dataa(\u1_m0_wo0_mtree_add0_4_o[11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_2_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_2_o[10]~38 ),
	.combout(\u1_m0_wo0_mtree_add1_2_o[11]~39_combout ),
	.cout(\u1_m0_wo0_mtree_add1_2_o[11]~40 ));
defparam \u1_m0_wo0_mtree_add1_2_o[11]~39 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_2_o[11]~39 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_2_o[12]~41 (
	.dataa(\u1_m0_wo0_mtree_add0_4_o[12]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_2_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_2_o[11]~40 ),
	.combout(\u1_m0_wo0_mtree_add1_2_o[12]~41_combout ),
	.cout(\u1_m0_wo0_mtree_add1_2_o[12]~42 ));
defparam \u1_m0_wo0_mtree_add1_2_o[12]~41 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_2_o[12]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_2_o[13]~43 (
	.dataa(\u1_m0_wo0_mtree_add0_4_o[13]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_2_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_2_o[12]~42 ),
	.combout(\u1_m0_wo0_mtree_add1_2_o[13]~43_combout ),
	.cout(\u1_m0_wo0_mtree_add1_2_o[13]~44 ));
defparam \u1_m0_wo0_mtree_add1_2_o[13]~43 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_2_o[13]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_2_o[14]~45 (
	.dataa(\u1_m0_wo0_mtree_add0_4_o[14]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_2_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_2_o[13]~44 ),
	.combout(\u1_m0_wo0_mtree_add1_2_o[14]~45_combout ),
	.cout(\u1_m0_wo0_mtree_add1_2_o[14]~46 ));
defparam \u1_m0_wo0_mtree_add1_2_o[14]~45 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_2_o[14]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_2_o[15]~47 (
	.dataa(\u1_m0_wo0_mtree_add0_4_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_2_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_2_o[14]~46 ),
	.combout(\u1_m0_wo0_mtree_add1_2_o[15]~47_combout ),
	.cout(\u1_m0_wo0_mtree_add1_2_o[15]~48 ));
defparam \u1_m0_wo0_mtree_add1_2_o[15]~47 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_2_o[15]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_2_o[17]~49 (
	.dataa(\u1_m0_wo0_mtree_add0_4_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_10_sub_2_o[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_add1_2_o[15]~48 ),
	.combout(\u1_m0_wo0_mtree_add1_2_o[17]~49_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_add1_2_o[17]~49 .lut_mask = 16'h6969;
defparam \u1_m0_wo0_mtree_add1_2_o[17]~49 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add1_2_o[17] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_2_o[17]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_2_o[17]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_2_o[17] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_2_o[17] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_1_o[10]~31 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][10]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_1_o[9]~30 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_1_o[10]~31_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_1_o[10]~32 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[10]~31 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[10]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_1_o[11]~33 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][10]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_1_o[10]~32 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_1_o[11]~33_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_1_o[11]~34 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[11]~33 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[11]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_1_o[12]~35 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr18|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_1_o[11]~34 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_1_o[12]~35_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_1_o[12]~36 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[12]~35 .lut_mask = 16'hF0AA;
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[12]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_1_o[13]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_1_o[12]~36 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_1_o[13]~37_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[13]~37 .lut_mask = 16'hF0F0;
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[13]~37 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_12_add_1_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_1_o[13]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_1_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_1_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_1_o[12]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_1_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_1_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_1_o[11]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_1_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_1_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_1_o[10]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_1_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_3_o[10]~27 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][7]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_12_add_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_3_o[9]~26 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_3_o[10]~27_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_3_o[10]~28 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[10]~27 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[10]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_3_o[11]~29 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][8]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_12_add_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_3_o[10]~28 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_3_o[11]~29_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_3_o[11]~30 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[11]~29 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[11]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_3_o[12]~31 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][9]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_12_add_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_3_o[11]~30 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_3_o[12]~31_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_3_o[12]~32 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[12]~31 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[12]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_3_o[13]~33 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][10]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_12_add_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_3_o[12]~32 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_3_o[13]~33_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_3_o[13]~34 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[13]~33 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[13]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_3_o[14]~35 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_12_add_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_3_o[13]~34 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_3_o[14]~35_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_12_add_3_o[14]~36 ));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[14]~35 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[14]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_12_add_3_o[15]~37 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr18_q_11|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_12_add_1_o[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_12_add_3_o[14]~36 ),
	.combout(\u1_m0_wo0_mtree_mult1_12_add_3_o[15]~37_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[15]~37 .lut_mask = 16'h6969;
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[15]~37 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_12_add_3_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_3_o[15]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_3_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[15] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_1_o[10]~33 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][7]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_1_o[9]~32 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[10]~33_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[10]~34 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[10]~33 .lut_mask = 16'h694D;
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[10]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_1_o[11]~35 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][8]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_1_o[10]~34 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[11]~35_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[11]~36 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[11]~35 .lut_mask = 16'h962B;
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[11]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_1_o[12]~37 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][9]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_1_o[11]~36 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[12]~37_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[12]~38 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[12]~37 .lut_mask = 16'h694D;
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[12]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_1_o[13]~39 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][10]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr17|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_1_o[12]~38 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[13]~39_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[13]~40 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[13]~39 .lut_mask = 16'h962B;
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[13]~39 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_1_o[14]~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_1_o[13]~40 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[14]~41_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[14]~42 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[14]~41 .lut_mask = 16'h0F0F;
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[14]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_1_o[15]~43 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_1_o[14]~42 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_1_o[15]~43_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[15]~43 .lut_mask = 16'hF0F0;
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[15]~43 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_1_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[15]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_1_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_1_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[14]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_1_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_1_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[13]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_1_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_1_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[12]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_1_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_1_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[11]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_1_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_1_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_1_o[10]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_1_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_3_o[10]~23 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][5]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_3_o[9]~22 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[10]~23_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[10]~24 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[10]~23 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[10]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_3_o[11]~25 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][6]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_3_o[10]~24 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[11]~25_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[11]~26 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[11]~25 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[11]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_3_o[12]~27 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][7]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_3_o[11]~26 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[12]~27_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[12]~28 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[12]~27 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[12]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_3_o[13]~29 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][8]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_3_o[12]~28 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[13]~29_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[13]~30 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[13]~29 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[13]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_3_o[14]~31 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][9]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_3_o[13]~30 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[14]~31_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[14]~32 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[14]~31 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[14]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_3_o[15]~33 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][10]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_1_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_3_o[14]~32 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[15]~33_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[15]~34 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[15]~33 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[15]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_3_o[16]~35 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_1_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_3_o[15]~34 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[16]~35_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[16]~36 ));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[16]~35 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[16]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_13_sub_3_o[17]~37 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr17_q_11|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_1_o[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_13_sub_3_o[16]~36 ),
	.combout(\u1_m0_wo0_mtree_mult1_13_sub_3_o[17]~37_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[17]~37 .lut_mask = 16'h9696;
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[17]~37 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_3_o[17] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_3_o[17]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_3_o[17]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[17] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[17] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_3_o[16] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_3_o[16]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_3_o[16]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[16] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[16] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_3_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_3_o[15]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_3_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_3_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_3_o[14]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_3_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_3_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_3_o[14]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_3_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_3_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_3_o[13]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_3_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_3_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_3_o[13]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_3_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_3_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_3_o[12]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_3_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_3_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_3_o[12]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_3_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_3_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_3_o[11]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_3_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_3_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_3_o[11]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_3_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_12_add_3_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_12_add_3_o[10]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_12_add_3_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_12_add_3_o[10] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_13_sub_3_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_13_sub_3_o[10]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_13_sub_3_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_13_sub_3_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_6_o[10]~39 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_3_o[10]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_3_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_6_o[9]~38 ),
	.combout(\u1_m0_wo0_mtree_add0_6_o[10]~39_combout ),
	.cout(\u1_m0_wo0_mtree_add0_6_o[10]~40 ));
defparam \u1_m0_wo0_mtree_add0_6_o[10]~39 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_6_o[10]~39 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_6_o[11]~41 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_3_o[11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_3_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_6_o[10]~40 ),
	.combout(\u1_m0_wo0_mtree_add0_6_o[11]~41_combout ),
	.cout(\u1_m0_wo0_mtree_add0_6_o[11]~42 ));
defparam \u1_m0_wo0_mtree_add0_6_o[11]~41 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_6_o[11]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_6_o[12]~43 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_3_o[12]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_3_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_6_o[11]~42 ),
	.combout(\u1_m0_wo0_mtree_add0_6_o[12]~43_combout ),
	.cout(\u1_m0_wo0_mtree_add0_6_o[12]~44 ));
defparam \u1_m0_wo0_mtree_add0_6_o[12]~43 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_6_o[12]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_6_o[13]~45 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_3_o[13]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_3_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_6_o[12]~44 ),
	.combout(\u1_m0_wo0_mtree_add0_6_o[13]~45_combout ),
	.cout(\u1_m0_wo0_mtree_add0_6_o[13]~46 ));
defparam \u1_m0_wo0_mtree_add0_6_o[13]~45 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_6_o[13]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_6_o[14]~47 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_3_o[14]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_3_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_6_o[13]~46 ),
	.combout(\u1_m0_wo0_mtree_add0_6_o[14]~47_combout ),
	.cout(\u1_m0_wo0_mtree_add0_6_o[14]~48 ));
defparam \u1_m0_wo0_mtree_add0_6_o[14]~47 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_6_o[14]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_6_o[15]~49 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_3_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_3_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_6_o[14]~48 ),
	.combout(\u1_m0_wo0_mtree_add0_6_o[15]~49_combout ),
	.cout(\u1_m0_wo0_mtree_add0_6_o[15]~50 ));
defparam \u1_m0_wo0_mtree_add0_6_o[15]~49 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_6_o[15]~49 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_6_o[16]~51 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_3_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_3_o[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_6_o[15]~50 ),
	.combout(\u1_m0_wo0_mtree_add0_6_o[16]~51_combout ),
	.cout(\u1_m0_wo0_mtree_add0_6_o[16]~52 ));
defparam \u1_m0_wo0_mtree_add0_6_o[16]~51 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_6_o[16]~51 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_6_o[17]~53 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_3_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_3_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_6_o[16]~52 ),
	.combout(\u1_m0_wo0_mtree_add0_6_o[17]~53_combout ),
	.cout(\u1_m0_wo0_mtree_add0_6_o[17]~54 ));
defparam \u1_m0_wo0_mtree_add0_6_o[17]~53 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_6_o[17]~53 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_6_o[18]~55 (
	.dataa(\u1_m0_wo0_mtree_mult1_12_add_3_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_13_sub_3_o[17]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_add0_6_o[17]~54 ),
	.combout(\u1_m0_wo0_mtree_add0_6_o[18]~55_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_add0_6_o[18]~55 .lut_mask = 16'h6969;
defparam \u1_m0_wo0_mtree_add0_6_o[18]~55 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add0_6_o[18] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_6_o[18]~55_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_6_o[18]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_6_o[18] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_6_o[18] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_1_o[10]~29 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][8]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_1_o[9]~28 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_1_o[10]~29_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_1_o[10]~30 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[10]~29 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[10]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_1_o[11]~31 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][9]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_1_o[10]~30 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_1_o[11]~31_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_1_o[11]~32 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[11]~31 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[11]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_1_o[12]~33 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][10]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_1_o[11]~32 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_1_o[12]~33_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_1_o[12]~34 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[12]~33 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[12]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_1_o[13]~35 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr16|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_1_o[12]~34 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_1_o[13]~35_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_1_o[13]~36 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[13]~35 .lut_mask = 16'hF0AA;
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[13]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_1_o[14]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_1_o[13]~36 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_1_o[14]~37_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[14]~37 .lut_mask = 16'hF0F0;
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[14]~37 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_14_add_1_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_1_o[14]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_1_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_1_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_1_o[13]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_1_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_1_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_1_o[12]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_1_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_1_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_1_o[11]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_1_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_1_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_1_o[10]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_1_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_3_o[10]~23 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][5]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_14_add_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_3_o[9]~22 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_3_o[10]~23_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_3_o[10]~24 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[10]~23 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[10]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_3_o[11]~25 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][6]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_14_add_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_3_o[10]~24 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_3_o[11]~25_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_3_o[11]~26 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[11]~25 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[11]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_3_o[12]~27 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][7]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_14_add_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_3_o[11]~26 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_3_o[12]~27_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_3_o[12]~28 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[12]~27 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[12]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_3_o[13]~29 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][8]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_14_add_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_3_o[12]~28 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_3_o[13]~29_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_3_o[13]~30 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[13]~29 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[13]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_3_o[14]~31 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][9]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_14_add_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_3_o[13]~30 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_3_o[14]~31_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_3_o[14]~32 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[14]~31 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[14]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_3_o[15]~33 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][10]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_14_add_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_3_o[14]~32 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_3_o[15]~33_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_3_o[15]~34 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[15]~33 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[15]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_3_o[16]~35 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_14_add_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_3_o[15]~34 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_3_o[16]~35_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_14_add_3_o[16]~36 ));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[16]~35 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[16]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_14_add_3_o[17]~37 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr16_q_11|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_14_add_1_o[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_14_add_3_o[16]~36 ),
	.combout(\u1_m0_wo0_mtree_mult1_14_add_3_o[17]~37_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[17]~37 .lut_mask = 16'h6969;
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[17]~37 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_14_add_3_o[17] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_3_o[17]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_3_o[17]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[17] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[17] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_15_sub_1_o[10]~37 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][3]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_15_sub_1_o[9]~36 ),
	.combout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[10]~37_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[10]~38 ));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[10]~37 .lut_mask = 16'h694D;
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[10]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_15_sub_1_o[11]~39 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][4]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_15_sub_1_o[10]~38 ),
	.combout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[11]~39_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[11]~40 ));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[11]~39 .lut_mask = 16'h962B;
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[11]~39 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_15_sub_1_o[12]~41 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][5]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_15_sub_1_o[11]~40 ),
	.combout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[12]~41_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[12]~42 ));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[12]~41 .lut_mask = 16'h694D;
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[12]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_15_sub_1_o[13]~43 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][6]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_15_sub_1_o[12]~42 ),
	.combout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[13]~43_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[13]~44 ));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[13]~43 .lut_mask = 16'h962B;
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[13]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_15_sub_1_o[14]~45 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][7]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_15_sub_1_o[13]~44 ),
	.combout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[14]~45_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[14]~46 ));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[14]~45 .lut_mask = 16'h694D;
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[14]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_15_sub_1_o[15]~47 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][8]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_15_sub_1_o[14]~46 ),
	.combout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[15]~47_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[15]~48 ));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[15]~47 .lut_mask = 16'h962B;
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[15]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_15_sub_1_o[16]~49 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][9]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_15_sub_1_o[15]~48 ),
	.combout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[16]~49_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[16]~50 ));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[16]~49 .lut_mask = 16'h694D;
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[16]~49 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_15_sub_1_o[17]~51 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][10]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr15_q_11|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_15_sub_1_o[16]~50 ),
	.combout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[17]~51_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[17]~52 ));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[17]~51 .lut_mask = 16'h962B;
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[17]~51 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_15_sub_1_o[18]~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_15_sub_1_o[17]~52 ),
	.combout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[18]~53_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[18]~54 ));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[18]~53 .lut_mask = 16'h0F0F;
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[18]~53 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_15_sub_1_o[19]~55 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_15_sub_1_o[18]~54 ),
	.combout(\u1_m0_wo0_mtree_mult1_15_sub_1_o[19]~55_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[19]~55 .lut_mask = 16'hF0F0;
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[19]~55 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[19] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_15_sub_1_o[19]~55_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[19]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[19] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[19] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[18] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_15_sub_1_o[18]~53_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[18]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[18] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[18] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[17] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_15_sub_1_o[17]~51_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[17]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[17] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[17] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_3_o[16] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_3_o[16]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_3_o[16]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[16] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[16] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[16] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_15_sub_1_o[16]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[16]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[16] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[16] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_3_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_3_o[15]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_3_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_15_sub_1_o[15]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_3_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_3_o[14]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_3_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_15_sub_1_o[14]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_3_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_3_o[13]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_3_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_15_sub_1_o[13]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_3_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_3_o[12]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_3_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_15_sub_1_o[12]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_3_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_3_o[11]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_3_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_15_sub_1_o[11]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_14_add_3_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_14_add_3_o[10]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_14_add_3_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_14_add_3_o[10] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_15_sub_1_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_15_sub_1_o[10]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_15_sub_1_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_15_sub_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[10]~41 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[10]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_7_o[9]~40 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[10]~41_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[10]~42 ));
defparam \u1_m0_wo0_mtree_add0_7_o[10]~41 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_7_o[10]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[11]~43 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_7_o[10]~42 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[11]~43_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[11]~44 ));
defparam \u1_m0_wo0_mtree_add0_7_o[11]~43 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_7_o[11]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[12]~45 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[12]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_7_o[11]~44 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[12]~45_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[12]~46 ));
defparam \u1_m0_wo0_mtree_add0_7_o[12]~45 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_7_o[12]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[13]~47 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[13]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_7_o[12]~46 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[13]~47_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[13]~48 ));
defparam \u1_m0_wo0_mtree_add0_7_o[13]~47 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_7_o[13]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[14]~49 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[14]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_7_o[13]~48 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[14]~49_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[14]~50 ));
defparam \u1_m0_wo0_mtree_add0_7_o[14]~49 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_7_o[14]~49 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[15]~51 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_7_o[14]~50 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[15]~51_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[15]~52 ));
defparam \u1_m0_wo0_mtree_add0_7_o[15]~51 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_7_o[15]~51 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[16]~53 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[16]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_7_o[15]~52 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[16]~53_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[16]~54 ));
defparam \u1_m0_wo0_mtree_add0_7_o[16]~53 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_7_o[16]~53 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[17]~55 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[17]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_7_o[16]~54 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[17]~55_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[17]~56 ));
defparam \u1_m0_wo0_mtree_add0_7_o[17]~55 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_7_o[17]~55 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[18]~57 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[17]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[18]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_7_o[17]~56 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[18]~57_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[18]~58 ));
defparam \u1_m0_wo0_mtree_add0_7_o[18]~57 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_7_o[18]~57 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[19]~59 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[17]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[19]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_7_o[18]~58 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[19]~59_combout ),
	.cout(\u1_m0_wo0_mtree_add0_7_o[19]~60 ));
defparam \u1_m0_wo0_mtree_add0_7_o[19]~59 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_7_o[19]~59 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_7_o[20]~61 (
	.dataa(\u1_m0_wo0_mtree_mult1_14_add_3_o[17]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_15_sub_1_o[19]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_add0_7_o[19]~60 ),
	.combout(\u1_m0_wo0_mtree_add0_7_o[20]~61_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_add0_7_o[20]~61 .lut_mask = 16'h6969;
defparam \u1_m0_wo0_mtree_add0_7_o[20]~61 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add0_7_o[20] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[20]~61_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[20]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[20] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[20] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_7_o[19] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[19]~59_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[19]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[19] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[19] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_7_o[18] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[18]~57_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[18]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[18] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[18] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_6_o[17] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_6_o[17]~53_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_6_o[17]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_6_o[17] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_6_o[17] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_7_o[17] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[17]~55_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[17]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[17] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[17] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_6_o[16] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_6_o[16]~51_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_6_o[16]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_6_o[16] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_6_o[16] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_7_o[16] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[16]~53_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[16]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[16] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[16] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_6_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_6_o[15]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_6_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_6_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_6_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_7_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[15]~51_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_6_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_6_o[14]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_6_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_6_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_6_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_7_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[14]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_6_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_6_o[13]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_6_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_6_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_6_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_7_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[13]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_6_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_6_o[12]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_6_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_6_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_6_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_7_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[12]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_6_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_6_o[11]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_6_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_6_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_6_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_7_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[11]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_6_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_6_o[10]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_6_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_6_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_6_o[10] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_7_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_7_o[10]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_7_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_7_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_7_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[10]~41 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[10]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_3_o[9]~40 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[10]~41_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[10]~42 ));
defparam \u1_m0_wo0_mtree_add1_3_o[10]~41 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_3_o[10]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[11]~43 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[11]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_3_o[10]~42 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[11]~43_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[11]~44 ));
defparam \u1_m0_wo0_mtree_add1_3_o[11]~43 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_3_o[11]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[12]~45 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[12]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_3_o[11]~44 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[12]~45_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[12]~46 ));
defparam \u1_m0_wo0_mtree_add1_3_o[12]~45 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_3_o[12]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[13]~47 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[13]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_3_o[12]~46 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[13]~47_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[13]~48 ));
defparam \u1_m0_wo0_mtree_add1_3_o[13]~47 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_3_o[13]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[14]~49 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[14]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_3_o[13]~48 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[14]~49_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[14]~50 ));
defparam \u1_m0_wo0_mtree_add1_3_o[14]~49 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_3_o[14]~49 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[15]~51 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_3_o[14]~50 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[15]~51_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[15]~52 ));
defparam \u1_m0_wo0_mtree_add1_3_o[15]~51 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_3_o[15]~51 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[16]~53 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[16]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_3_o[15]~52 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[16]~53_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[16]~54 ));
defparam \u1_m0_wo0_mtree_add1_3_o[16]~53 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_3_o[16]~53 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[17]~55 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[17]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_3_o[16]~54 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[17]~55_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[17]~56 ));
defparam \u1_m0_wo0_mtree_add1_3_o[17]~55 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_3_o[17]~55 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[18]~57 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[18]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[18]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_3_o[17]~56 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[18]~57_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[18]~58 ));
defparam \u1_m0_wo0_mtree_add1_3_o[18]~57 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_3_o[18]~57 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[19]~59 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[18]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[19]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_3_o[18]~58 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[19]~59_combout ),
	.cout(\u1_m0_wo0_mtree_add1_3_o[19]~60 ));
defparam \u1_m0_wo0_mtree_add1_3_o[19]~59 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_3_o[19]~59 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_3_o[20]~61 (
	.dataa(\u1_m0_wo0_mtree_add0_6_o[18]~q ),
	.datab(\u1_m0_wo0_mtree_add0_7_o[20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_add1_3_o[19]~60 ),
	.combout(\u1_m0_wo0_mtree_add1_3_o[20]~61_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_add1_3_o[20]~61 .lut_mask = 16'h6969;
defparam \u1_m0_wo0_mtree_add1_3_o[20]~61 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add1_3_o[20] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[20]~61_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[20]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[20] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[20] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_3_o[19] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[19]~59_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[19]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[19] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[19] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_3_o[18] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[18]~57_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[18]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[18] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[18] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_3_o[17] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[17]~55_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[17]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[17] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[17] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_3_o[16] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[16]~53_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[16]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[16] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[16] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_2_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_2_o[15]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_2_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_2_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_2_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_3_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[15]~51_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_2_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_2_o[14]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_2_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_2_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_2_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_3_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[14]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_2_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_2_o[13]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_2_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_2_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_2_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_3_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[13]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_2_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_2_o[12]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_2_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_2_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_2_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_3_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[12]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_2_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_2_o[11]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_2_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_2_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_2_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_3_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[11]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_2_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_2_o[10]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_2_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_2_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_2_o[10] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_3_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_3_o[10]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_3_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_3_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_3_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[10]~41 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[10]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_1_o[9]~40 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[10]~41_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[10]~42 ));
defparam \u1_m0_wo0_mtree_add2_1_o[10]~41 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add2_1_o[10]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[11]~43 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[11]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_1_o[10]~42 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[11]~43_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[11]~44 ));
defparam \u1_m0_wo0_mtree_add2_1_o[11]~43 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_1_o[11]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[12]~45 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[12]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_1_o[11]~44 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[12]~45_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[12]~46 ));
defparam \u1_m0_wo0_mtree_add2_1_o[12]~45 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add2_1_o[12]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[13]~47 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[13]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_1_o[12]~46 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[13]~47_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[13]~48 ));
defparam \u1_m0_wo0_mtree_add2_1_o[13]~47 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_1_o[13]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[14]~49 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[14]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_1_o[13]~48 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[14]~49_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[14]~50 ));
defparam \u1_m0_wo0_mtree_add2_1_o[14]~49 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add2_1_o[14]~49 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[15]~51 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_1_o[14]~50 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[15]~51_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[15]~52 ));
defparam \u1_m0_wo0_mtree_add2_1_o[15]~51 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_1_o[15]~51 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[16]~53 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[17]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_1_o[15]~52 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[16]~53_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[16]~54 ));
defparam \u1_m0_wo0_mtree_add2_1_o[16]~53 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add2_1_o[16]~53 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[17]~55 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[17]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_1_o[16]~54 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[17]~55_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[17]~56 ));
defparam \u1_m0_wo0_mtree_add2_1_o[17]~55 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_1_o[17]~55 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[18]~57 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[17]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[18]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_1_o[17]~56 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[18]~57_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[18]~58 ));
defparam \u1_m0_wo0_mtree_add2_1_o[18]~57 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add2_1_o[18]~57 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[19]~59 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[17]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[19]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_1_o[18]~58 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[19]~59_combout ),
	.cout(\u1_m0_wo0_mtree_add2_1_o[19]~60 ));
defparam \u1_m0_wo0_mtree_add2_1_o[19]~59 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_1_o[19]~59 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_1_o[20]~61 (
	.dataa(\u1_m0_wo0_mtree_add1_2_o[17]~q ),
	.datab(\u1_m0_wo0_mtree_add1_3_o[20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_add2_1_o[19]~60 ),
	.combout(\u1_m0_wo0_mtree_add2_1_o[20]~61_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_add2_1_o[20]~61 .lut_mask = 16'h6969;
defparam \u1_m0_wo0_mtree_add2_1_o[20]~61 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add2_1_o[20] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[20]~61_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[20]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[20] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[20] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_1_o[19] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[19]~59_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[19]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[19] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[19] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_1_o[18] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[18]~57_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[18]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[18] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[18] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_1_o[17] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[17]~55_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[17]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[17] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[17] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_1_o[16] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[16]~53_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[16]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[16] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[16] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_1_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[15]~51_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_1_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[14]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_1_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[13]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_1_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_1_o[12]~38_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_1_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_1_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_1_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_1_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[12]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_1_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_1_o[11]~36_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_1_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_1_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_1_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_1_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[11]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_1_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_1_o[10]~34_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_1_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_1_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_1_o[10] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_1_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_1_o[10]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_1_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_1_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[10]~41 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[10]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_0_o[9]~40 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[10]~41_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[10]~42 ));
defparam \u1_m0_wo0_mtree_add3_0_o[10]~41 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add3_0_o[10]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[11]~43 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[11]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_0_o[10]~42 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[11]~43_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[11]~44 ));
defparam \u1_m0_wo0_mtree_add3_0_o[11]~43 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_0_o[11]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[12]~45 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[12]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_0_o[11]~44 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[12]~45_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[12]~46 ));
defparam \u1_m0_wo0_mtree_add3_0_o[12]~45 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add3_0_o[12]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[13]~47 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_0_o[12]~46 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[13]~47_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[13]~48 ));
defparam \u1_m0_wo0_mtree_add3_0_o[13]~47 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_0_o[13]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[14]~49 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_0_o[13]~48 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[14]~49_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[14]~50 ));
defparam \u1_m0_wo0_mtree_add3_0_o[14]~49 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add3_0_o[14]~49 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[15]~51 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_0_o[14]~50 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[15]~51_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[15]~52 ));
defparam \u1_m0_wo0_mtree_add3_0_o[15]~51 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_0_o[15]~51 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[16]~53 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_0_o[15]~52 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[16]~53_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[16]~54 ));
defparam \u1_m0_wo0_mtree_add3_0_o[16]~53 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add3_0_o[16]~53 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[17]~55 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_0_o[16]~54 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[17]~55_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[17]~56 ));
defparam \u1_m0_wo0_mtree_add3_0_o[17]~55 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_0_o[17]~55 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[18]~57 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[18]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_0_o[17]~56 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[18]~57_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[18]~58 ));
defparam \u1_m0_wo0_mtree_add3_0_o[18]~57 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add3_0_o[18]~57 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[19]~59 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[19]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_0_o[18]~58 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[19]~59_combout ),
	.cout(\u1_m0_wo0_mtree_add3_0_o[19]~60 ));
defparam \u1_m0_wo0_mtree_add3_0_o[19]~59 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_0_o[19]~59 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_0_o[20]~61 (
	.dataa(\u1_m0_wo0_mtree_add1_1_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_add2_1_o[20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_add3_0_o[19]~60 ),
	.combout(\u1_m0_wo0_mtree_add3_0_o[20]~61_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_add3_0_o[20]~61 .lut_mask = 16'h6969;
defparam \u1_m0_wo0_mtree_add3_0_o[20]~61 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add3_0_o[20] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[20]~61_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[20]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[20] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[20] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_1_o[10]~29 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][8]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_1_o[9]~28 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_1_o[10]~29_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_1_o[10]~30 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[10]~29 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[10]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_1_o[11]~31 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][9]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_1_o[10]~30 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_1_o[11]~31_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_1_o[11]~32 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[11]~31 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[11]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_1_o[12]~33 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][10]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_1_o[11]~32 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_1_o[12]~33_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_1_o[12]~34 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[12]~33 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[12]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_1_o[13]~35 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr14|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_1_o[12]~34 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_1_o[13]~35_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_1_o[13]~36 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[13]~35 .lut_mask = 16'hF0AA;
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[13]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_1_o[14]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_1_o[13]~36 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_1_o[14]~37_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[14]~37 .lut_mask = 16'hF0F0;
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[14]~37 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_16_add_1_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_1_o[14]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_1_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_1_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_1_o[13]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_1_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_1_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_1_o[12]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_1_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_1_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_1_o[11]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_1_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_1_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_1_o[10]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_1_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_3_o[10]~23 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][5]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_16_add_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_3_o[9]~22 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_3_o[10]~23_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_3_o[10]~24 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[10]~23 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[10]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_3_o[11]~25 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][6]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_16_add_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_3_o[10]~24 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_3_o[11]~25_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_3_o[11]~26 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[11]~25 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[11]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_3_o[12]~27 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][7]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_16_add_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_3_o[11]~26 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_3_o[12]~27_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_3_o[12]~28 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[12]~27 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[12]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_3_o[13]~29 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][8]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_16_add_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_3_o[12]~28 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_3_o[13]~29_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_3_o[13]~30 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[13]~29 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[13]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_3_o[14]~31 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][9]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_16_add_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_3_o[13]~30 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_3_o[14]~31_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_3_o[14]~32 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[14]~31 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[14]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_3_o[15]~33 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][10]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_16_add_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_3_o[14]~32 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_3_o[15]~33_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_3_o[15]~34 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[15]~33 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[15]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_3_o[16]~35 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_16_add_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_3_o[15]~34 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_3_o[16]~35_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_16_add_3_o[16]~36 ));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[16]~35 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[16]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_16_add_3_o[17]~37 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr14_q_11|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_16_add_1_o[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_16_add_3_o[16]~36 ),
	.combout(\u1_m0_wo0_mtree_mult1_16_add_3_o[17]~37_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[17]~37 .lut_mask = 16'h6969;
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[17]~37 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_16_add_3_o[17] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_3_o[17]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_3_o[17]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[17] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[17] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_1_o[10]~33 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][7]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_1_o[9]~32 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[10]~33_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[10]~34 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[10]~33 .lut_mask = 16'h694D;
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[10]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_1_o[11]~35 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][8]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_1_o[10]~34 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[11]~35_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[11]~36 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[11]~35 .lut_mask = 16'h962B;
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[11]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_1_o[12]~37 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][9]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_1_o[11]~36 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[12]~37_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[12]~38 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[12]~37 .lut_mask = 16'h694D;
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[12]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_1_o[13]~39 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][10]~q ),
	.datab(\u1_m0_wo0_wi0_r0_delayr13|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_1_o[12]~38 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[13]~39_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[13]~40 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[13]~39 .lut_mask = 16'h962B;
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[13]~39 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_1_o[14]~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_1_o[13]~40 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[14]~41_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[14]~42 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[14]~41 .lut_mask = 16'h0F0F;
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[14]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_1_o[15]~43 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_1_o[14]~42 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_1_o[15]~43_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[15]~43 .lut_mask = 16'hF0F0;
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[15]~43 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_1_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[15]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_1_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_1_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[14]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_1_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_1_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[13]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_1_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_1_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[12]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_1_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_1_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[11]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_1_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_1_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_1_o[10]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_1_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_3_o[10]~23 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][5]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_3_o[9]~22 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[10]~23_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[10]~24 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[10]~23 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[10]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_3_o[11]~25 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][6]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_3_o[10]~24 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[11]~25_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[11]~26 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[11]~25 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[11]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_3_o[12]~27 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][7]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_3_o[11]~26 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[12]~27_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[12]~28 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[12]~27 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[12]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_3_o[13]~29 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][8]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_3_o[12]~28 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[13]~29_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[13]~30 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[13]~29 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[13]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_3_o[14]~31 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][9]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_3_o[13]~30 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[14]~31_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[14]~32 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[14]~31 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[14]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_3_o[15]~33 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][10]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_1_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_3_o[14]~32 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[15]~33_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[15]~34 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[15]~33 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[15]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_3_o[16]~35 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_1_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_3_o[15]~34 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[16]~35_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[16]~36 ));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[16]~35 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[16]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_17_sub_3_o[17]~37 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr13_q_11|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_1_o[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_17_sub_3_o[16]~36 ),
	.combout(\u1_m0_wo0_mtree_mult1_17_sub_3_o[17]~37_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[17]~37 .lut_mask = 16'h9696;
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[17]~37 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_3_o[17] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_3_o[17]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_3_o[17]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[17] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[17] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_3_o[16] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_3_o[16]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_3_o[16]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[16] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[16] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_3_o[16] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_3_o[16]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_3_o[16]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[16] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[16] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_3_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_3_o[15]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_3_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_3_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_3_o[15]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_3_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_3_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_3_o[14]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_3_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_3_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_3_o[14]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_3_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_3_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_3_o[13]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_3_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_3_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_3_o[13]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_3_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_3_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_3_o[12]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_3_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_3_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_3_o[12]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_3_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_3_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_3_o[11]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_3_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_3_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_3_o[11]~25_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_3_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_16_add_3_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_16_add_3_o[10]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_16_add_3_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_16_add_3_o[10] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_17_sub_3_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_17_sub_3_o[10]~23_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_17_sub_3_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_17_sub_3_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_8_o[10]~39 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_3_o[10]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_3_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_8_o[9]~38 ),
	.combout(\u1_m0_wo0_mtree_add0_8_o[10]~39_combout ),
	.cout(\u1_m0_wo0_mtree_add0_8_o[10]~40 ));
defparam \u1_m0_wo0_mtree_add0_8_o[10]~39 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_8_o[10]~39 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_8_o[11]~41 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_3_o[11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_3_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_8_o[10]~40 ),
	.combout(\u1_m0_wo0_mtree_add0_8_o[11]~41_combout ),
	.cout(\u1_m0_wo0_mtree_add0_8_o[11]~42 ));
defparam \u1_m0_wo0_mtree_add0_8_o[11]~41 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_8_o[11]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_8_o[12]~43 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_3_o[12]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_3_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_8_o[11]~42 ),
	.combout(\u1_m0_wo0_mtree_add0_8_o[12]~43_combout ),
	.cout(\u1_m0_wo0_mtree_add0_8_o[12]~44 ));
defparam \u1_m0_wo0_mtree_add0_8_o[12]~43 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_8_o[12]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_8_o[13]~45 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_3_o[13]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_3_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_8_o[12]~44 ),
	.combout(\u1_m0_wo0_mtree_add0_8_o[13]~45_combout ),
	.cout(\u1_m0_wo0_mtree_add0_8_o[13]~46 ));
defparam \u1_m0_wo0_mtree_add0_8_o[13]~45 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_8_o[13]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_8_o[14]~47 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_3_o[14]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_3_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_8_o[13]~46 ),
	.combout(\u1_m0_wo0_mtree_add0_8_o[14]~47_combout ),
	.cout(\u1_m0_wo0_mtree_add0_8_o[14]~48 ));
defparam \u1_m0_wo0_mtree_add0_8_o[14]~47 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_8_o[14]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_8_o[15]~49 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_3_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_3_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_8_o[14]~48 ),
	.combout(\u1_m0_wo0_mtree_add0_8_o[15]~49_combout ),
	.cout(\u1_m0_wo0_mtree_add0_8_o[15]~50 ));
defparam \u1_m0_wo0_mtree_add0_8_o[15]~49 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_8_o[15]~49 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_8_o[16]~51 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_3_o[16]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_3_o[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_8_o[15]~50 ),
	.combout(\u1_m0_wo0_mtree_add0_8_o[16]~51_combout ),
	.cout(\u1_m0_wo0_mtree_add0_8_o[16]~52 ));
defparam \u1_m0_wo0_mtree_add0_8_o[16]~51 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_8_o[16]~51 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_8_o[17]~53 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_3_o[17]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_3_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_8_o[16]~52 ),
	.combout(\u1_m0_wo0_mtree_add0_8_o[17]~53_combout ),
	.cout(\u1_m0_wo0_mtree_add0_8_o[17]~54 ));
defparam \u1_m0_wo0_mtree_add0_8_o[17]~53 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_8_o[17]~53 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_8_o[18]~55 (
	.dataa(\u1_m0_wo0_mtree_mult1_16_add_3_o[17]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_17_sub_3_o[17]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_add0_8_o[17]~54 ),
	.combout(\u1_m0_wo0_mtree_add0_8_o[18]~55_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_add0_8_o[18]~55 .lut_mask = 16'h6969;
defparam \u1_m0_wo0_mtree_add0_8_o[18]~55 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add0_8_o[18] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_8_o[18]~55_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_8_o[18]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_8_o[18] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_8_o[18] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_1_o[10]~31 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][10]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_1_o[9]~30 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_1_o[10]~31_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_1_o[10]~32 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[10]~31 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[10]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_1_o[11]~33 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][10]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_1_o[10]~32 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_1_o[11]~33_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_1_o[11]~34 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[11]~33 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[11]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_1_o[12]~35 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_11|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_1_o[11]~34 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_1_o[12]~35_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_1_o[12]~36 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[12]~35 .lut_mask = 16'hF0AA;
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[12]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_1_o[13]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_1_o[12]~36 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_1_o[13]~37_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[13]~37 .lut_mask = 16'hF0F0;
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[13]~37 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_18_add_1_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_1_o[13]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_1_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_1_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_1_o[12]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_1_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_1_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_1_o[11]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_1_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_1_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_1_o[10]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_1_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_3_o[10]~27 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][7]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_3_o[9]~26 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_3_o[10]~27_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_3_o[10]~28 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[10]~27 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[10]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_3_o[11]~29 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][8]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_3_o[10]~28 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_3_o[11]~29_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_3_o[11]~30 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[11]~29 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[11]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_3_o[12]~31 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][9]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_3_o[11]~30 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_3_o[12]~31_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_3_o[12]~32 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[12]~31 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[12]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_3_o[13]~33 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][10]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_3_o[12]~32 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_3_o[13]~33_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_3_o[13]~34 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[13]~33 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[13]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_3_o[14]~35 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_3_o[13]~34 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_3_o[14]~35_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_18_add_3_o[14]~36 ));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[14]~35 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[14]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_18_add_3_o[15]~37 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr12_q_12|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_1_o[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_18_add_3_o[14]~36 ),
	.combout(\u1_m0_wo0_mtree_mult1_18_add_3_o[15]~37_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[15]~37 .lut_mask = 16'h6969;
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[15]~37 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_18_add_3_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_3_o[15]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_3_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_8_o[17] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_8_o[17]~53_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_8_o[17]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_8_o[17] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_8_o[17] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_8_o[16] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_8_o[16]~51_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_8_o[16]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_8_o[16] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_8_o[16] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_8_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_8_o[15]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_8_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_8_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_8_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_8_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_8_o[14]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_8_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_8_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_8_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_3_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_3_o[14]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_3_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_8_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_8_o[13]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_8_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_8_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_8_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_3_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_3_o[13]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_3_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_8_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_8_o[12]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_8_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_8_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_8_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_3_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_3_o[12]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_3_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_8_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_8_o[11]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_8_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_8_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_8_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_3_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_3_o[11]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_3_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_8_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_8_o[10]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_8_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_8_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_8_o[10] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_18_add_3_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_18_add_3_o[10]~27_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_18_add_3_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_18_add_3_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[10]~40 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[10]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_4_o[9]~39 ),
	.combout(\u1_m0_wo0_mtree_add1_4_o[10]~40_combout ),
	.cout(\u1_m0_wo0_mtree_add1_4_o[10]~41 ));
defparam \u1_m0_wo0_mtree_add1_4_o[10]~40 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_4_o[10]~40 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[11]~42 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_4_o[10]~41 ),
	.combout(\u1_m0_wo0_mtree_add1_4_o[11]~42_combout ),
	.cout(\u1_m0_wo0_mtree_add1_4_o[11]~43 ));
defparam \u1_m0_wo0_mtree_add1_4_o[11]~42 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_4_o[11]~42 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[12]~44 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[12]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_4_o[11]~43 ),
	.combout(\u1_m0_wo0_mtree_add1_4_o[12]~44_combout ),
	.cout(\u1_m0_wo0_mtree_add1_4_o[12]~45 ));
defparam \u1_m0_wo0_mtree_add1_4_o[12]~44 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_4_o[12]~44 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[13]~46 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[13]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_4_o[12]~45 ),
	.combout(\u1_m0_wo0_mtree_add1_4_o[13]~46_combout ),
	.cout(\u1_m0_wo0_mtree_add1_4_o[13]~47 ));
defparam \u1_m0_wo0_mtree_add1_4_o[13]~46 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_4_o[13]~46 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[14]~48 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[14]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_4_o[13]~47 ),
	.combout(\u1_m0_wo0_mtree_add1_4_o[14]~48_combout ),
	.cout(\u1_m0_wo0_mtree_add1_4_o[14]~49 ));
defparam \u1_m0_wo0_mtree_add1_4_o[14]~48 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_4_o[14]~48 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[15]~50 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_4_o[14]~49 ),
	.combout(\u1_m0_wo0_mtree_add1_4_o[15]~50_combout ),
	.cout(\u1_m0_wo0_mtree_add1_4_o[15]~51 ));
defparam \u1_m0_wo0_mtree_add1_4_o[15]~50 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_4_o[15]~50 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[16]~52 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[16]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_4_o[15]~51 ),
	.combout(\u1_m0_wo0_mtree_add1_4_o[16]~52_combout ),
	.cout(\u1_m0_wo0_mtree_add1_4_o[16]~53 ));
defparam \u1_m0_wo0_mtree_add1_4_o[16]~52 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_4_o[16]~52 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[17]~54 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[17]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_4_o[16]~53 ),
	.combout(\u1_m0_wo0_mtree_add1_4_o[17]~54_combout ),
	.cout(\u1_m0_wo0_mtree_add1_4_o[17]~55 ));
defparam \u1_m0_wo0_mtree_add1_4_o[17]~54 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_4_o[17]~54 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[18]~56 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[18]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_4_o[17]~55 ),
	.combout(\u1_m0_wo0_mtree_add1_4_o[18]~56_combout ),
	.cout(\u1_m0_wo0_mtree_add1_4_o[18]~57 ));
defparam \u1_m0_wo0_mtree_add1_4_o[18]~56 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_4_o[18]~56 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_4_o[20]~58 (
	.dataa(\u1_m0_wo0_mtree_add0_8_o[18]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_18_add_3_o[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_add1_4_o[18]~57 ),
	.combout(\u1_m0_wo0_mtree_add1_4_o[20]~58_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_add1_4_o[20]~58 .lut_mask = 16'h9696;
defparam \u1_m0_wo0_mtree_add1_4_o[20]~58 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add1_4_o[20] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[20]~58_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[20]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[20] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[20] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_0_o[10]~30 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_0_o[9]~29 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[10]~30_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[10]~31 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[10]~30 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[10]~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_0_o[11]~32 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_0_o[10]~31 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[11]~32_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[11]~33 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[11]~32 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[11]~32 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_0_o[12]~34 (
	.dataa(\u1_m0_wo0_wi0_r0_delayr10|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_0_o[11]~33 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_0_o[12]~34_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[12]~34 .lut_mask = 16'hA5A5;
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[12]~34 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_0_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_0_o[12]~34_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_0_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_0_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_0_o[11]~32_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_0_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_0_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_0_o[10]~30_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_0_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_0_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_2_o[10]~29 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][8]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_20_sub_0_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_2_o[9]~28 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[10]~29_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[10]~30 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[10]~29 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[10]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_2_o[11]~31 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][9]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_20_sub_0_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_2_o[10]~30 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[11]~31_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[11]~32 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[11]~31 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[11]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_2_o[12]~33 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][10]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_20_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_2_o[11]~32 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[12]~33_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[12]~34 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[12]~33 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[12]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_2_o[13]~35 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_20_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_2_o[12]~34 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[13]~35_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[13]~36 ));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[13]~35 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[13]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_20_sub_2_o[14]~37 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr10_q_11|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_20_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_20_sub_2_o[13]~36 ),
	.combout(\u1_m0_wo0_mtree_mult1_20_sub_2_o[14]~37_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[14]~37 .lut_mask = 16'h9696;
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[14]~37 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_2_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_2_o[14]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_2_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[14] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_21_add_1_o[9]~29 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][8]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_21_add_1_o[8]~28 ),
	.combout(\u1_m0_wo0_mtree_mult1_21_add_1_o[9]~29_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_21_add_1_o[9]~30 ));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[9]~29 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[9]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_21_add_1_o[10]~31 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][10]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_21_add_1_o[9]~30 ),
	.combout(\u1_m0_wo0_mtree_mult1_21_add_1_o[10]~31_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_21_add_1_o[10]~32 ));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[10]~31 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[10]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_21_add_1_o[11]~33 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][10]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_21_add_1_o[10]~32 ),
	.combout(\u1_m0_wo0_mtree_mult1_21_add_1_o[11]~33_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_21_add_1_o[11]~34 ));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[11]~33 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[11]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_21_add_1_o[12]~35 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr9_q_11|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_21_add_1_o[11]~34 ),
	.combout(\u1_m0_wo0_mtree_mult1_21_add_1_o[12]~35_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_21_add_1_o[12]~36 ));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[12]~35 .lut_mask = 16'hF0AA;
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[12]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_21_add_1_o[13]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_21_add_1_o[12]~36 ),
	.combout(\u1_m0_wo0_mtree_mult1_21_add_1_o[13]~37_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[13]~37 .lut_mask = 16'hF0F0;
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[13]~37 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_21_add_1_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_21_add_1_o[13]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_21_add_1_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_2_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_2_o[13]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_2_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_21_add_1_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_21_add_1_o[12]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_21_add_1_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_2_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_2_o[12]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_2_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_21_add_1_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_21_add_1_o[11]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_21_add_1_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_2_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_2_o[11]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_2_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_21_add_1_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_21_add_1_o[10]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_21_add_1_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[10] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_20_sub_2_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_20_sub_2_o[10]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_20_sub_2_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_20_sub_2_o[10] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_21_add_1_o[9] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_21_add_1_o[9]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_21_add_1_o[9]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[9] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_21_add_1_o[9] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_10_o[10]~33 (
	.dataa(\u1_m0_wo0_mtree_mult1_20_sub_2_o[10]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_21_add_1_o[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_10_o[9]~32 ),
	.combout(\u1_m0_wo0_mtree_add0_10_o[10]~33_combout ),
	.cout(\u1_m0_wo0_mtree_add0_10_o[10]~34 ));
defparam \u1_m0_wo0_mtree_add0_10_o[10]~33 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_10_o[10]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_10_o[11]~35 (
	.dataa(\u1_m0_wo0_mtree_mult1_20_sub_2_o[11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_21_add_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_10_o[10]~34 ),
	.combout(\u1_m0_wo0_mtree_add0_10_o[11]~35_combout ),
	.cout(\u1_m0_wo0_mtree_add0_10_o[11]~36 ));
defparam \u1_m0_wo0_mtree_add0_10_o[11]~35 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_10_o[11]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_10_o[12]~37 (
	.dataa(\u1_m0_wo0_mtree_mult1_20_sub_2_o[12]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_21_add_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_10_o[11]~36 ),
	.combout(\u1_m0_wo0_mtree_add0_10_o[12]~37_combout ),
	.cout(\u1_m0_wo0_mtree_add0_10_o[12]~38 ));
defparam \u1_m0_wo0_mtree_add0_10_o[12]~37 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_10_o[12]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_10_o[13]~39 (
	.dataa(\u1_m0_wo0_mtree_mult1_20_sub_2_o[13]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_21_add_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_10_o[12]~38 ),
	.combout(\u1_m0_wo0_mtree_add0_10_o[13]~39_combout ),
	.cout(\u1_m0_wo0_mtree_add0_10_o[13]~40 ));
defparam \u1_m0_wo0_mtree_add0_10_o[13]~39 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_10_o[13]~39 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_10_o[14]~41 (
	.dataa(\u1_m0_wo0_mtree_mult1_20_sub_2_o[14]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_21_add_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_10_o[13]~40 ),
	.combout(\u1_m0_wo0_mtree_add0_10_o[14]~41_combout ),
	.cout(\u1_m0_wo0_mtree_add0_10_o[14]~42 ));
defparam \u1_m0_wo0_mtree_add0_10_o[14]~41 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_10_o[14]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_10_o[15]~43 (
	.dataa(\u1_m0_wo0_mtree_mult1_20_sub_2_o[14]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_21_add_1_o[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_add0_10_o[14]~42 ),
	.combout(\u1_m0_wo0_mtree_add0_10_o[15]~43_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_add0_10_o[15]~43 .lut_mask = 16'h6969;
defparam \u1_m0_wo0_mtree_add0_10_o[15]~43 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add0_10_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_10_o[15]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_10_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_10_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_10_o[15] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_22_sub_1_o[10]~29 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][8]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_22_sub_1_o[9]~28 ),
	.combout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[10]~29_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[10]~30 ));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[10]~29 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[10]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_22_sub_1_o[11]~31 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][9]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_22_sub_1_o[10]~30 ),
	.combout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[11]~31_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[11]~32 ));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[11]~31 .lut_mask = 16'h692B;
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[11]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_22_sub_1_o[12]~33 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][10]~q ),
	.datab(\d_u1_m0_wo0_wi0_r0_delayr8_q_12|delay_signals[0][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_22_sub_1_o[11]~32 ),
	.combout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[12]~33_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[12]~34 ));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[12]~33 .lut_mask = 16'h964D;
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[12]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_22_sub_1_o[13]~35 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_22_sub_1_o[12]~34 ),
	.combout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[13]~35_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[13]~36 ));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[13]~35 .lut_mask = 16'h0F0F;
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[13]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_22_sub_1_o[14]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_22_sub_1_o[13]~36 ),
	.combout(\u1_m0_wo0_mtree_mult1_22_sub_1_o[14]~37_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[14]~37 .lut_mask = 16'hF0F0;
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[14]~37 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_22_sub_1_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_22_sub_1_o[14]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_22_sub_1_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_10_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_10_o[14]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_10_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_10_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_10_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_10_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_10_o[13]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_10_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_10_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_10_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_22_sub_1_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_22_sub_1_o[13]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_22_sub_1_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_10_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_10_o[12]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_10_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_10_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_10_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_22_sub_1_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_22_sub_1_o[12]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_22_sub_1_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_10_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_10_o[11]~35_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_10_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_10_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_10_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_22_sub_1_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_22_sub_1_o[11]~31_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_22_sub_1_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_10_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_10_o[10]~33_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_10_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_10_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_10_o[10] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_22_sub_1_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_22_sub_1_o[10]~29_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_22_sub_1_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_22_sub_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_5_o[10]~37 (
	.dataa(\u1_m0_wo0_mtree_add0_10_o[10]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_22_sub_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_5_o[9]~36 ),
	.combout(\u1_m0_wo0_mtree_add1_5_o[10]~37_combout ),
	.cout(\u1_m0_wo0_mtree_add1_5_o[10]~38 ));
defparam \u1_m0_wo0_mtree_add1_5_o[10]~37 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_5_o[10]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_5_o[11]~39 (
	.dataa(\u1_m0_wo0_mtree_add0_10_o[11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_22_sub_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_5_o[10]~38 ),
	.combout(\u1_m0_wo0_mtree_add1_5_o[11]~39_combout ),
	.cout(\u1_m0_wo0_mtree_add1_5_o[11]~40 ));
defparam \u1_m0_wo0_mtree_add1_5_o[11]~39 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_5_o[11]~39 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_5_o[12]~41 (
	.dataa(\u1_m0_wo0_mtree_add0_10_o[12]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_22_sub_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_5_o[11]~40 ),
	.combout(\u1_m0_wo0_mtree_add1_5_o[12]~41_combout ),
	.cout(\u1_m0_wo0_mtree_add1_5_o[12]~42 ));
defparam \u1_m0_wo0_mtree_add1_5_o[12]~41 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_5_o[12]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_5_o[13]~43 (
	.dataa(\u1_m0_wo0_mtree_add0_10_o[13]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_22_sub_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_5_o[12]~42 ),
	.combout(\u1_m0_wo0_mtree_add1_5_o[13]~43_combout ),
	.cout(\u1_m0_wo0_mtree_add1_5_o[13]~44 ));
defparam \u1_m0_wo0_mtree_add1_5_o[13]~43 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_5_o[13]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_5_o[14]~45 (
	.dataa(\u1_m0_wo0_mtree_add0_10_o[14]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_22_sub_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_5_o[13]~44 ),
	.combout(\u1_m0_wo0_mtree_add1_5_o[14]~45_combout ),
	.cout(\u1_m0_wo0_mtree_add1_5_o[14]~46 ));
defparam \u1_m0_wo0_mtree_add1_5_o[14]~45 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add1_5_o[14]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_5_o[15]~47 (
	.dataa(\u1_m0_wo0_mtree_add0_10_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_22_sub_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add1_5_o[14]~46 ),
	.combout(\u1_m0_wo0_mtree_add1_5_o[15]~47_combout ),
	.cout(\u1_m0_wo0_mtree_add1_5_o[15]~48 ));
defparam \u1_m0_wo0_mtree_add1_5_o[15]~47 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add1_5_o[15]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add1_5_o[17]~49 (
	.dataa(\u1_m0_wo0_mtree_add0_10_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_22_sub_1_o[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_add1_5_o[15]~48 ),
	.combout(\u1_m0_wo0_mtree_add1_5_o[17]~49_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_add1_5_o[17]~49 .lut_mask = 16'h6969;
defparam \u1_m0_wo0_mtree_add1_5_o[17]~49 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add1_5_o[17] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_5_o[17]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_5_o[17]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_5_o[17] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_5_o[17] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_4_o[18] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[18]~56_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[18]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[18] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[18] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_4_o[17] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[17]~54_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[17]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[17] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[17] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_4_o[16] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[16]~52_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[16]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[16] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[16] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_4_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[15]~50_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_5_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_5_o[15]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_5_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_5_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_5_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_4_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[14]~48_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_5_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_5_o[14]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_5_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_5_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_5_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_4_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[13]~46_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_5_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_5_o[13]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_5_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_5_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_5_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_4_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[12]~44_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_5_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_5_o[12]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_5_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_5_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_5_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_4_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[11]~42_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_5_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_5_o[11]~39_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_5_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_5_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_5_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_4_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_4_o[10]~40_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_4_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_4_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_4_o[10] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add1_5_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add1_5_o[10]~37_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add1_5_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add1_5_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add1_5_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[10]~41 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[10]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_2_o[9]~40 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[10]~41_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[10]~42 ));
defparam \u1_m0_wo0_mtree_add2_2_o[10]~41 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add2_2_o[10]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[11]~43 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[11]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_2_o[10]~42 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[11]~43_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[11]~44 ));
defparam \u1_m0_wo0_mtree_add2_2_o[11]~43 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_2_o[11]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[12]~45 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[12]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_2_o[11]~44 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[12]~45_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[12]~46 ));
defparam \u1_m0_wo0_mtree_add2_2_o[12]~45 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add2_2_o[12]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[13]~47 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[13]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_2_o[12]~46 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[13]~47_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[13]~48 ));
defparam \u1_m0_wo0_mtree_add2_2_o[13]~47 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_2_o[13]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[14]~49 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[14]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_2_o[13]~48 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[14]~49_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[14]~50 ));
defparam \u1_m0_wo0_mtree_add2_2_o[14]~49 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add2_2_o[14]~49 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[15]~51 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_2_o[14]~50 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[15]~51_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[15]~52 ));
defparam \u1_m0_wo0_mtree_add2_2_o[15]~51 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_2_o[15]~51 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[16]~53 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[16]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_2_o[15]~52 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[16]~53_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[16]~54 ));
defparam \u1_m0_wo0_mtree_add2_2_o[16]~53 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add2_2_o[16]~53 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[17]~55 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[17]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_2_o[16]~54 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[17]~55_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[17]~56 ));
defparam \u1_m0_wo0_mtree_add2_2_o[17]~55 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_2_o[17]~55 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[18]~57 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[18]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_2_o[17]~56 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[18]~57_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[18]~58 ));
defparam \u1_m0_wo0_mtree_add2_2_o[18]~57 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add2_2_o[18]~57 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[19]~59 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[20]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add2_2_o[18]~58 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[19]~59_combout ),
	.cout(\u1_m0_wo0_mtree_add2_2_o[19]~60 ));
defparam \u1_m0_wo0_mtree_add2_2_o[19]~59 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add2_2_o[19]~59 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add2_2_o[20]~61 (
	.dataa(\u1_m0_wo0_mtree_add1_4_o[20]~q ),
	.datab(\u1_m0_wo0_mtree_add1_5_o[17]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_add2_2_o[19]~60 ),
	.combout(\u1_m0_wo0_mtree_add2_2_o[20]~61_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_add2_2_o[20]~61 .lut_mask = 16'h6969;
defparam \u1_m0_wo0_mtree_add2_2_o[20]~61 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add2_2_o[20] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[20]~61_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[20]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[20] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[20] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_25_sub_0_o[10]~30 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_25_sub_0_o[9]~29 ),
	.combout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[10]~30_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[10]~31 ));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[10]~30 .lut_mask = 16'hA5AF;
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[10]~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_25_sub_0_o[11]~32 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_mult1_25_sub_0_o[10]~31 ),
	.combout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[11]~32_combout ),
	.cout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[11]~33 ));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[11]~32 .lut_mask = 16'h5A05;
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[11]~32 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_mult1_25_sub_0_o[12]~34 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr5_q_13|delay_signals[0][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_mult1_25_sub_0_o[11]~33 ),
	.combout(\u1_m0_wo0_mtree_mult1_25_sub_0_o[12]~34_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[12]~34 .lut_mask = 16'hA5A5;
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[12]~34 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_mult1_25_sub_0_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_25_sub_0_o[12]~34_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_25_sub_0_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_25_sub_0_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_25_sub_0_o[11]~32_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_25_sub_0_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_mult1_25_sub_0_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_mult1_25_sub_0_o[10]~30_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_mult1_25_sub_0_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_mult1_25_sub_0_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_12_o[10]~34 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][10]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_25_sub_0_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_12_o[9]~33 ),
	.combout(\u1_m0_wo0_mtree_add0_12_o[10]~34_combout ),
	.cout(\u1_m0_wo0_mtree_add0_12_o[10]~35 ));
defparam \u1_m0_wo0_mtree_add0_12_o[10]~34 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_12_o[10]~34 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_12_o[11]~36 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_25_sub_0_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_12_o[10]~35 ),
	.combout(\u1_m0_wo0_mtree_add0_12_o[11]~36_combout ),
	.cout(\u1_m0_wo0_mtree_add0_12_o[11]~37 ));
defparam \u1_m0_wo0_mtree_add0_12_o[11]~36 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add0_12_o[11]~36 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_12_o[12]~38 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_25_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add0_12_o[11]~37 ),
	.combout(\u1_m0_wo0_mtree_add0_12_o[12]~38_combout ),
	.cout(\u1_m0_wo0_mtree_add0_12_o[12]~39 ));
defparam \u1_m0_wo0_mtree_add0_12_o[12]~38 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add0_12_o[12]~38 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add0_12_o[13]~40 (
	.dataa(\d_u1_m0_wo0_wi0_r0_delayr6_q_14|delay_signals[0][11]~q ),
	.datab(\u1_m0_wo0_mtree_mult1_25_sub_0_o[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_add0_12_o[12]~39 ),
	.combout(\u1_m0_wo0_mtree_add0_12_o[13]~40_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_add0_12_o[13]~40 .lut_mask = 16'h9696;
defparam \u1_m0_wo0_mtree_add0_12_o[13]~40 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add0_12_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_12_o[13]~40_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_12_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_12_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_12_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_2_o[19] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[19]~59_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[19]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[19] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[19] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_2_o[18] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[18]~57_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[18]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[18] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[18] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_2_o[17] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[17]~55_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[17]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[17] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[17] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_2_o[16] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[16]~53_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[16]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[16] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[16] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_2_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[15]~51_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_2_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[14]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_2_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[13]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_2_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[12]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_12_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_12_o[12]~38_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_12_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_12_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_12_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_2_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[11]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_12_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_12_o[11]~36_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_12_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_12_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_12_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add2_2_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add2_2_o[10]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add2_2_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add2_2_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add2_2_o[10] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add0_12_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add0_12_o[10]~34_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add0_12_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add0_12_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add0_12_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[10]~41 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[10]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_1_o[9]~40 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[10]~41_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[10]~42 ));
defparam \u1_m0_wo0_mtree_add3_1_o[10]~41 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add3_1_o[10]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[11]~43 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[11]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_1_o[10]~42 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[11]~43_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[11]~44 ));
defparam \u1_m0_wo0_mtree_add3_1_o[11]~43 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_1_o[11]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[12]~45 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[12]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_1_o[11]~44 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[12]~45_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[12]~46 ));
defparam \u1_m0_wo0_mtree_add3_1_o[12]~45 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add3_1_o[12]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[13]~47 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[13]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_1_o[12]~46 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[13]~47_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[13]~48 ));
defparam \u1_m0_wo0_mtree_add3_1_o[13]~47 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_1_o[13]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[14]~49 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[14]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_1_o[13]~48 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[14]~49_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[14]~50 ));
defparam \u1_m0_wo0_mtree_add3_1_o[14]~49 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add3_1_o[14]~49 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[15]~51 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_1_o[14]~50 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[15]~51_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[15]~52 ));
defparam \u1_m0_wo0_mtree_add3_1_o[15]~51 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_1_o[15]~51 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[16]~53 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[16]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_1_o[15]~52 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[16]~53_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[16]~54 ));
defparam \u1_m0_wo0_mtree_add3_1_o[16]~53 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add3_1_o[16]~53 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[17]~55 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[17]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_1_o[16]~54 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[17]~55_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[17]~56 ));
defparam \u1_m0_wo0_mtree_add3_1_o[17]~55 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_1_o[17]~55 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[18]~57 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[18]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_1_o[17]~56 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[18]~57_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[18]~58 ));
defparam \u1_m0_wo0_mtree_add3_1_o[18]~57 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add3_1_o[18]~57 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[19]~59 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[19]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add3_1_o[18]~58 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[19]~59_combout ),
	.cout(\u1_m0_wo0_mtree_add3_1_o[19]~60 ));
defparam \u1_m0_wo0_mtree_add3_1_o[19]~59 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add3_1_o[19]~59 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add3_1_o[20]~61 (
	.dataa(\u1_m0_wo0_mtree_add2_2_o[20]~q ),
	.datab(\u1_m0_wo0_mtree_add0_12_o[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_add3_1_o[19]~60 ),
	.combout(\u1_m0_wo0_mtree_add3_1_o[20]~61_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_add3_1_o[20]~61 .lut_mask = 16'h6969;
defparam \u1_m0_wo0_mtree_add3_1_o[20]~61 .sum_lutc_input = "cin";

dffeas \u1_m0_wo0_mtree_add3_1_o[20] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[20]~61_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[20]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[20] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[20] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_0_o[19] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[19]~59_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[19]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[19] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[19] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_1_o[19] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[19]~59_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[19]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[19] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[19] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_0_o[18] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[18]~57_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[18]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[18] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[18] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_1_o[18] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[18]~57_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[18]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[18] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[18] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_0_o[17] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[17]~55_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[17]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[17] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[17] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_1_o[17] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[17]~55_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[17]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[17] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[17] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_0_o[16] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[16]~53_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[16]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[16] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[16] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_1_o[16] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[16]~53_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[16]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[16] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[16] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_0_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[15]~51_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_1_o[15] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[15]~51_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[15]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[15] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[15] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_0_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[14]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_1_o[14] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[14]~49_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[14]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[14] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[14] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_0_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[13]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_1_o[13] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[13]~47_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[13]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[13] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[13] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_0_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[12]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_1_o[12] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[12]~45_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[12]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[12] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[12] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_0_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[11]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_1_o[11] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[11]~43_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[11]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[11] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[11] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_0_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_0_o[10]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_0_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_0_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_0_o[10] .power_up = "low";

dffeas \u1_m0_wo0_mtree_add3_1_o[10] (
	.clk(clk),
	.d(\u1_m0_wo0_mtree_add3_1_o[10]~41_combout ),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\u1_m0_wo0_mtree_add3_1_o[10]~q ),
	.prn(vcc));
defparam \u1_m0_wo0_mtree_add3_1_o[10] .is_wysiwyg = "true";
defparam \u1_m0_wo0_mtree_add3_1_o[10] .power_up = "low";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[10]~32 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[10]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add4_0_o[9]~31 ),
	.combout(\u1_m0_wo0_mtree_add4_0_o[10]~32_combout ),
	.cout(\u1_m0_wo0_mtree_add4_0_o[10]~33 ));
defparam \u1_m0_wo0_mtree_add4_0_o[10]~32 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add4_0_o[10]~32 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[11]~34 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[11]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add4_0_o[10]~33 ),
	.combout(\u1_m0_wo0_mtree_add4_0_o[11]~34_combout ),
	.cout(\u1_m0_wo0_mtree_add4_0_o[11]~35 ));
defparam \u1_m0_wo0_mtree_add4_0_o[11]~34 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add4_0_o[11]~34 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[12]~36 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[12]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add4_0_o[11]~35 ),
	.combout(\u1_m0_wo0_mtree_add4_0_o[12]~36_combout ),
	.cout(\u1_m0_wo0_mtree_add4_0_o[12]~37 ));
defparam \u1_m0_wo0_mtree_add4_0_o[12]~36 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add4_0_o[12]~36 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[13]~38 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[13]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add4_0_o[12]~37 ),
	.combout(\u1_m0_wo0_mtree_add4_0_o[13]~38_combout ),
	.cout(\u1_m0_wo0_mtree_add4_0_o[13]~39 ));
defparam \u1_m0_wo0_mtree_add4_0_o[13]~38 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add4_0_o[13]~38 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[14]~40 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[14]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add4_0_o[13]~39 ),
	.combout(\u1_m0_wo0_mtree_add4_0_o[14]~40_combout ),
	.cout(\u1_m0_wo0_mtree_add4_0_o[14]~41 ));
defparam \u1_m0_wo0_mtree_add4_0_o[14]~40 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add4_0_o[14]~40 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[15]~42 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[15]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add4_0_o[14]~41 ),
	.combout(\u1_m0_wo0_mtree_add4_0_o[15]~42_combout ),
	.cout(\u1_m0_wo0_mtree_add4_0_o[15]~43 ));
defparam \u1_m0_wo0_mtree_add4_0_o[15]~42 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add4_0_o[15]~42 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[16]~44 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[16]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add4_0_o[15]~43 ),
	.combout(\u1_m0_wo0_mtree_add4_0_o[16]~44_combout ),
	.cout(\u1_m0_wo0_mtree_add4_0_o[16]~45 ));
defparam \u1_m0_wo0_mtree_add4_0_o[16]~44 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add4_0_o[16]~44 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[17]~46 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[17]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add4_0_o[16]~45 ),
	.combout(\u1_m0_wo0_mtree_add4_0_o[17]~46_combout ),
	.cout(\u1_m0_wo0_mtree_add4_0_o[17]~47 ));
defparam \u1_m0_wo0_mtree_add4_0_o[17]~46 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add4_0_o[17]~46 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[18]~48 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[18]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[18]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add4_0_o[17]~47 ),
	.combout(\u1_m0_wo0_mtree_add4_0_o[18]~48_combout ),
	.cout(\u1_m0_wo0_mtree_add4_0_o[18]~49 ));
defparam \u1_m0_wo0_mtree_add4_0_o[18]~48 .lut_mask = 16'h698E;
defparam \u1_m0_wo0_mtree_add4_0_o[18]~48 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[19]~50 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[19]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[19]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\u1_m0_wo0_mtree_add4_0_o[18]~49 ),
	.combout(\u1_m0_wo0_mtree_add4_0_o[19]~50_combout ),
	.cout(\u1_m0_wo0_mtree_add4_0_o[19]~51 ));
defparam \u1_m0_wo0_mtree_add4_0_o[19]~50 .lut_mask = 16'h9617;
defparam \u1_m0_wo0_mtree_add4_0_o[19]~50 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \u1_m0_wo0_mtree_add4_0_o[20]~52 (
	.dataa(\u1_m0_wo0_mtree_add3_0_o[20]~q ),
	.datab(\u1_m0_wo0_mtree_add3_1_o[20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\u1_m0_wo0_mtree_add4_0_o[19]~51 ),
	.combout(\u1_m0_wo0_mtree_add4_0_o[20]~52_combout ),
	.cout());
defparam \u1_m0_wo0_mtree_add4_0_o[20]~52 .lut_mask = 16'h6969;
defparam \u1_m0_wo0_mtree_add4_0_o[20]~52 .sum_lutc_input = "cin";

endmodule

module lms_dsp_dspba_delay (
	aclr,
	delay_signals_0_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_0_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_1 (
	aclr,
	delay_signals_0_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_0_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \delay_signals[1][0]~q ;


dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(\delay_signals[1][0]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[1][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][0]~q ),
	.prn(vcc));
defparam \delay_signals[1][0] .is_wysiwyg = "true";
defparam \delay_signals[1][0] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_2 (
	aclr,
	delay_signals_0_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_0_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \delay_signals[2][0]~q ;
wire \delay_signals[1][0]~q ;


dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(\delay_signals[1][0]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[2][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][0]~q ),
	.prn(vcc));
defparam \delay_signals[2][0] .is_wysiwyg = "true";
defparam \delay_signals[2][0] .power_up = "low";

dffeas \delay_signals[1][0] (
	.clk(clk),
	.d(\delay_signals[2][0]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][0]~q ),
	.prn(vcc));
defparam \delay_signals[1][0] .is_wysiwyg = "true";
defparam \delay_signals[1][0] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_5 (
	aclr,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	delay_signals_8_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_6 (
	aclr,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_9_0,
	delay_signals_7_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_11_0,
	delay_signals_10_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_9_0;
output 	delay_signals_7_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_7 (
	aclr,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_8 (
	aclr,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_9 (
	aclr,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_10 (
	aclr,
	delay_signals_2_0,
	delay_signals_9_0,
	delay_signals_1_0,
	delay_signals_8_0,
	delay_signals_0_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_10_0,
	delay_signals_11_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_2_0;
output 	delay_signals_9_0;
output 	delay_signals_1_0;
output 	delay_signals_8_0;
output 	delay_signals_0_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_10_0;
output 	delay_signals_11_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_11 (
	aclr,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_12 (
	aclr,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_13 (
	aclr,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_14 (
	aclr,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	delay_signals_8_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_15 (
	aclr,
	u0_m0_wo0_mtree_mult1_8_sub_1_o_1,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	xin,
	delay_signals_11_0,
	delay_signals_10_0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	u0_m0_wo0_mtree_mult1_8_sub_1_o_1;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
input 	[11:0] xin;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \delay_signals[1][9]~q ;
wire \delay_signals[1][8]~q ;
wire \delay_signals[1][7]~q ;
wire \delay_signals[1][6]~q ;
wire \delay_signals[1][5]~q ;
wire \delay_signals[1][4]~q ;
wire \delay_signals[1][3]~q ;
wire \delay_signals[1][2]~q ;
wire \delay_signals[1][11]~q ;
wire \delay_signals[1][10]~q ;


dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(\delay_signals[1][9]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(\delay_signals[1][8]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(\delay_signals[1][7]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(\delay_signals[1][6]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(\delay_signals[1][5]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(\delay_signals[1][4]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(\delay_signals[1][3]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(\delay_signals[1][2]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(u0_m0_wo0_mtree_mult1_8_sub_1_o_1),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(\delay_signals[1][11]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(\delay_signals[1][10]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[1][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][9]~q ),
	.prn(vcc));
defparam \delay_signals[1][9] .is_wysiwyg = "true";
defparam \delay_signals[1][9] .power_up = "low";

dffeas \delay_signals[1][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][8]~q ),
	.prn(vcc));
defparam \delay_signals[1][8] .is_wysiwyg = "true";
defparam \delay_signals[1][8] .power_up = "low";

dffeas \delay_signals[1][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][7]~q ),
	.prn(vcc));
defparam \delay_signals[1][7] .is_wysiwyg = "true";
defparam \delay_signals[1][7] .power_up = "low";

dffeas \delay_signals[1][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][6]~q ),
	.prn(vcc));
defparam \delay_signals[1][6] .is_wysiwyg = "true";
defparam \delay_signals[1][6] .power_up = "low";

dffeas \delay_signals[1][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][5]~q ),
	.prn(vcc));
defparam \delay_signals[1][5] .is_wysiwyg = "true";
defparam \delay_signals[1][5] .power_up = "low";

dffeas \delay_signals[1][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][4]~q ),
	.prn(vcc));
defparam \delay_signals[1][4] .is_wysiwyg = "true";
defparam \delay_signals[1][4] .power_up = "low";

dffeas \delay_signals[1][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][3]~q ),
	.prn(vcc));
defparam \delay_signals[1][3] .is_wysiwyg = "true";
defparam \delay_signals[1][3] .power_up = "low";

dffeas \delay_signals[1][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][2]~q ),
	.prn(vcc));
defparam \delay_signals[1][2] .is_wysiwyg = "true";
defparam \delay_signals[1][2] .power_up = "low";

dffeas \delay_signals[1][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][11]~q ),
	.prn(vcc));
defparam \delay_signals[1][11] .is_wysiwyg = "true";
defparam \delay_signals[1][11] .power_up = "low";

dffeas \delay_signals[1][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][10]~q ),
	.prn(vcc));
defparam \delay_signals[1][10] .is_wysiwyg = "true";
defparam \delay_signals[1][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_16 (
	aclr,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_11_0,
	delay_signals_10_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_17 (
	aclr,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \delay_signals[2][9]~q ;
wire \delay_signals[1][9]~q ;
wire \delay_signals[2][8]~q ;
wire \delay_signals[1][8]~q ;
wire \delay_signals[2][7]~q ;
wire \delay_signals[1][7]~q ;
wire \delay_signals[2][6]~q ;
wire \delay_signals[1][6]~q ;
wire \delay_signals[2][5]~q ;
wire \delay_signals[1][5]~q ;
wire \delay_signals[2][4]~q ;
wire \delay_signals[1][4]~q ;
wire \delay_signals[2][3]~q ;
wire \delay_signals[1][3]~q ;
wire \delay_signals[2][2]~q ;
wire \delay_signals[1][2]~q ;
wire \delay_signals[2][0]~q ;
wire \delay_signals[1][0]~q ;
wire \delay_signals[2][1]~q ;
wire \delay_signals[1][1]~q ;
wire \delay_signals[2][11]~q ;
wire \delay_signals[1][11]~q ;
wire \delay_signals[2][10]~q ;
wire \delay_signals[1][10]~q ;


dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(\delay_signals[1][9]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(\delay_signals[1][8]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(\delay_signals[1][7]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(\delay_signals[1][6]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(\delay_signals[1][5]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(\delay_signals[1][4]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(\delay_signals[1][3]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(\delay_signals[1][2]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(\delay_signals[1][0]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(\delay_signals[1][1]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(\delay_signals[1][11]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(\delay_signals[1][10]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[2][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][9]~q ),
	.prn(vcc));
defparam \delay_signals[2][9] .is_wysiwyg = "true";
defparam \delay_signals[2][9] .power_up = "low";

dffeas \delay_signals[1][9] (
	.clk(clk),
	.d(\delay_signals[2][9]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][9]~q ),
	.prn(vcc));
defparam \delay_signals[1][9] .is_wysiwyg = "true";
defparam \delay_signals[1][9] .power_up = "low";

dffeas \delay_signals[2][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][8]~q ),
	.prn(vcc));
defparam \delay_signals[2][8] .is_wysiwyg = "true";
defparam \delay_signals[2][8] .power_up = "low";

dffeas \delay_signals[1][8] (
	.clk(clk),
	.d(\delay_signals[2][8]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][8]~q ),
	.prn(vcc));
defparam \delay_signals[1][8] .is_wysiwyg = "true";
defparam \delay_signals[1][8] .power_up = "low";

dffeas \delay_signals[2][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][7]~q ),
	.prn(vcc));
defparam \delay_signals[2][7] .is_wysiwyg = "true";
defparam \delay_signals[2][7] .power_up = "low";

dffeas \delay_signals[1][7] (
	.clk(clk),
	.d(\delay_signals[2][7]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][7]~q ),
	.prn(vcc));
defparam \delay_signals[1][7] .is_wysiwyg = "true";
defparam \delay_signals[1][7] .power_up = "low";

dffeas \delay_signals[2][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][6]~q ),
	.prn(vcc));
defparam \delay_signals[2][6] .is_wysiwyg = "true";
defparam \delay_signals[2][6] .power_up = "low";

dffeas \delay_signals[1][6] (
	.clk(clk),
	.d(\delay_signals[2][6]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][6]~q ),
	.prn(vcc));
defparam \delay_signals[1][6] .is_wysiwyg = "true";
defparam \delay_signals[1][6] .power_up = "low";

dffeas \delay_signals[2][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][5]~q ),
	.prn(vcc));
defparam \delay_signals[2][5] .is_wysiwyg = "true";
defparam \delay_signals[2][5] .power_up = "low";

dffeas \delay_signals[1][5] (
	.clk(clk),
	.d(\delay_signals[2][5]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][5]~q ),
	.prn(vcc));
defparam \delay_signals[1][5] .is_wysiwyg = "true";
defparam \delay_signals[1][5] .power_up = "low";

dffeas \delay_signals[2][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][4]~q ),
	.prn(vcc));
defparam \delay_signals[2][4] .is_wysiwyg = "true";
defparam \delay_signals[2][4] .power_up = "low";

dffeas \delay_signals[1][4] (
	.clk(clk),
	.d(\delay_signals[2][4]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][4]~q ),
	.prn(vcc));
defparam \delay_signals[1][4] .is_wysiwyg = "true";
defparam \delay_signals[1][4] .power_up = "low";

dffeas \delay_signals[2][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][3]~q ),
	.prn(vcc));
defparam \delay_signals[2][3] .is_wysiwyg = "true";
defparam \delay_signals[2][3] .power_up = "low";

dffeas \delay_signals[1][3] (
	.clk(clk),
	.d(\delay_signals[2][3]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][3]~q ),
	.prn(vcc));
defparam \delay_signals[1][3] .is_wysiwyg = "true";
defparam \delay_signals[1][3] .power_up = "low";

dffeas \delay_signals[2][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][2]~q ),
	.prn(vcc));
defparam \delay_signals[2][2] .is_wysiwyg = "true";
defparam \delay_signals[2][2] .power_up = "low";

dffeas \delay_signals[1][2] (
	.clk(clk),
	.d(\delay_signals[2][2]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][2]~q ),
	.prn(vcc));
defparam \delay_signals[1][2] .is_wysiwyg = "true";
defparam \delay_signals[1][2] .power_up = "low";

dffeas \delay_signals[2][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][0]~q ),
	.prn(vcc));
defparam \delay_signals[2][0] .is_wysiwyg = "true";
defparam \delay_signals[2][0] .power_up = "low";

dffeas \delay_signals[1][0] (
	.clk(clk),
	.d(\delay_signals[2][0]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][0]~q ),
	.prn(vcc));
defparam \delay_signals[1][0] .is_wysiwyg = "true";
defparam \delay_signals[1][0] .power_up = "low";

dffeas \delay_signals[2][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][1]~q ),
	.prn(vcc));
defparam \delay_signals[2][1] .is_wysiwyg = "true";
defparam \delay_signals[2][1] .power_up = "low";

dffeas \delay_signals[1][1] (
	.clk(clk),
	.d(\delay_signals[2][1]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][1]~q ),
	.prn(vcc));
defparam \delay_signals[1][1] .is_wysiwyg = "true";
defparam \delay_signals[1][1] .power_up = "low";

dffeas \delay_signals[2][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][11]~q ),
	.prn(vcc));
defparam \delay_signals[2][11] .is_wysiwyg = "true";
defparam \delay_signals[2][11] .power_up = "low";

dffeas \delay_signals[1][11] (
	.clk(clk),
	.d(\delay_signals[2][11]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][11]~q ),
	.prn(vcc));
defparam \delay_signals[1][11] .is_wysiwyg = "true";
defparam \delay_signals[1][11] .power_up = "low";

dffeas \delay_signals[2][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][10]~q ),
	.prn(vcc));
defparam \delay_signals[2][10] .is_wysiwyg = "true";
defparam \delay_signals[2][10] .power_up = "low";

dffeas \delay_signals[1][10] (
	.clk(clk),
	.d(\delay_signals[2][10]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][10]~q ),
	.prn(vcc));
defparam \delay_signals[1][10] .is_wysiwyg = "true";
defparam \delay_signals[1][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_18 (
	aclr,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_11_0,
	delay_signals_10_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \delay_signals[3][9]~q ;
wire \delay_signals[2][9]~q ;
wire \delay_signals[1][9]~q ;
wire \delay_signals[3][8]~q ;
wire \delay_signals[2][8]~q ;
wire \delay_signals[1][8]~q ;
wire \delay_signals[3][7]~q ;
wire \delay_signals[2][7]~q ;
wire \delay_signals[1][7]~q ;
wire \delay_signals[3][6]~q ;
wire \delay_signals[2][6]~q ;
wire \delay_signals[1][6]~q ;
wire \delay_signals[3][5]~q ;
wire \delay_signals[2][5]~q ;
wire \delay_signals[1][5]~q ;
wire \delay_signals[3][4]~q ;
wire \delay_signals[2][4]~q ;
wire \delay_signals[1][4]~q ;
wire \delay_signals[3][3]~q ;
wire \delay_signals[2][3]~q ;
wire \delay_signals[1][3]~q ;
wire \delay_signals[3][2]~q ;
wire \delay_signals[2][2]~q ;
wire \delay_signals[1][2]~q ;
wire \delay_signals[3][1]~q ;
wire \delay_signals[2][1]~q ;
wire \delay_signals[1][1]~q ;
wire \delay_signals[3][0]~q ;
wire \delay_signals[2][0]~q ;
wire \delay_signals[1][0]~q ;
wire \delay_signals[3][11]~q ;
wire \delay_signals[2][11]~q ;
wire \delay_signals[1][11]~q ;
wire \delay_signals[3][10]~q ;
wire \delay_signals[2][10]~q ;
wire \delay_signals[1][10]~q ;


dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(\delay_signals[1][9]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(\delay_signals[1][8]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(\delay_signals[1][7]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(\delay_signals[1][6]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(\delay_signals[1][5]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(\delay_signals[1][4]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(\delay_signals[1][3]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(\delay_signals[1][2]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(\delay_signals[1][1]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(\delay_signals[1][0]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(\delay_signals[1][11]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(\delay_signals[1][10]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[3][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][9]~q ),
	.prn(vcc));
defparam \delay_signals[3][9] .is_wysiwyg = "true";
defparam \delay_signals[3][9] .power_up = "low";

dffeas \delay_signals[2][9] (
	.clk(clk),
	.d(\delay_signals[3][9]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][9]~q ),
	.prn(vcc));
defparam \delay_signals[2][9] .is_wysiwyg = "true";
defparam \delay_signals[2][9] .power_up = "low";

dffeas \delay_signals[1][9] (
	.clk(clk),
	.d(\delay_signals[2][9]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][9]~q ),
	.prn(vcc));
defparam \delay_signals[1][9] .is_wysiwyg = "true";
defparam \delay_signals[1][9] .power_up = "low";

dffeas \delay_signals[3][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][8]~q ),
	.prn(vcc));
defparam \delay_signals[3][8] .is_wysiwyg = "true";
defparam \delay_signals[3][8] .power_up = "low";

dffeas \delay_signals[2][8] (
	.clk(clk),
	.d(\delay_signals[3][8]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][8]~q ),
	.prn(vcc));
defparam \delay_signals[2][8] .is_wysiwyg = "true";
defparam \delay_signals[2][8] .power_up = "low";

dffeas \delay_signals[1][8] (
	.clk(clk),
	.d(\delay_signals[2][8]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][8]~q ),
	.prn(vcc));
defparam \delay_signals[1][8] .is_wysiwyg = "true";
defparam \delay_signals[1][8] .power_up = "low";

dffeas \delay_signals[3][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][7]~q ),
	.prn(vcc));
defparam \delay_signals[3][7] .is_wysiwyg = "true";
defparam \delay_signals[3][7] .power_up = "low";

dffeas \delay_signals[2][7] (
	.clk(clk),
	.d(\delay_signals[3][7]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][7]~q ),
	.prn(vcc));
defparam \delay_signals[2][7] .is_wysiwyg = "true";
defparam \delay_signals[2][7] .power_up = "low";

dffeas \delay_signals[1][7] (
	.clk(clk),
	.d(\delay_signals[2][7]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][7]~q ),
	.prn(vcc));
defparam \delay_signals[1][7] .is_wysiwyg = "true";
defparam \delay_signals[1][7] .power_up = "low";

dffeas \delay_signals[3][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][6]~q ),
	.prn(vcc));
defparam \delay_signals[3][6] .is_wysiwyg = "true";
defparam \delay_signals[3][6] .power_up = "low";

dffeas \delay_signals[2][6] (
	.clk(clk),
	.d(\delay_signals[3][6]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][6]~q ),
	.prn(vcc));
defparam \delay_signals[2][6] .is_wysiwyg = "true";
defparam \delay_signals[2][6] .power_up = "low";

dffeas \delay_signals[1][6] (
	.clk(clk),
	.d(\delay_signals[2][6]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][6]~q ),
	.prn(vcc));
defparam \delay_signals[1][6] .is_wysiwyg = "true";
defparam \delay_signals[1][6] .power_up = "low";

dffeas \delay_signals[3][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][5]~q ),
	.prn(vcc));
defparam \delay_signals[3][5] .is_wysiwyg = "true";
defparam \delay_signals[3][5] .power_up = "low";

dffeas \delay_signals[2][5] (
	.clk(clk),
	.d(\delay_signals[3][5]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][5]~q ),
	.prn(vcc));
defparam \delay_signals[2][5] .is_wysiwyg = "true";
defparam \delay_signals[2][5] .power_up = "low";

dffeas \delay_signals[1][5] (
	.clk(clk),
	.d(\delay_signals[2][5]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][5]~q ),
	.prn(vcc));
defparam \delay_signals[1][5] .is_wysiwyg = "true";
defparam \delay_signals[1][5] .power_up = "low";

dffeas \delay_signals[3][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][4]~q ),
	.prn(vcc));
defparam \delay_signals[3][4] .is_wysiwyg = "true";
defparam \delay_signals[3][4] .power_up = "low";

dffeas \delay_signals[2][4] (
	.clk(clk),
	.d(\delay_signals[3][4]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][4]~q ),
	.prn(vcc));
defparam \delay_signals[2][4] .is_wysiwyg = "true";
defparam \delay_signals[2][4] .power_up = "low";

dffeas \delay_signals[1][4] (
	.clk(clk),
	.d(\delay_signals[2][4]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][4]~q ),
	.prn(vcc));
defparam \delay_signals[1][4] .is_wysiwyg = "true";
defparam \delay_signals[1][4] .power_up = "low";

dffeas \delay_signals[3][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][3]~q ),
	.prn(vcc));
defparam \delay_signals[3][3] .is_wysiwyg = "true";
defparam \delay_signals[3][3] .power_up = "low";

dffeas \delay_signals[2][3] (
	.clk(clk),
	.d(\delay_signals[3][3]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][3]~q ),
	.prn(vcc));
defparam \delay_signals[2][3] .is_wysiwyg = "true";
defparam \delay_signals[2][3] .power_up = "low";

dffeas \delay_signals[1][3] (
	.clk(clk),
	.d(\delay_signals[2][3]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][3]~q ),
	.prn(vcc));
defparam \delay_signals[1][3] .is_wysiwyg = "true";
defparam \delay_signals[1][3] .power_up = "low";

dffeas \delay_signals[3][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][2]~q ),
	.prn(vcc));
defparam \delay_signals[3][2] .is_wysiwyg = "true";
defparam \delay_signals[3][2] .power_up = "low";

dffeas \delay_signals[2][2] (
	.clk(clk),
	.d(\delay_signals[3][2]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][2]~q ),
	.prn(vcc));
defparam \delay_signals[2][2] .is_wysiwyg = "true";
defparam \delay_signals[2][2] .power_up = "low";

dffeas \delay_signals[1][2] (
	.clk(clk),
	.d(\delay_signals[2][2]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][2]~q ),
	.prn(vcc));
defparam \delay_signals[1][2] .is_wysiwyg = "true";
defparam \delay_signals[1][2] .power_up = "low";

dffeas \delay_signals[3][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][1]~q ),
	.prn(vcc));
defparam \delay_signals[3][1] .is_wysiwyg = "true";
defparam \delay_signals[3][1] .power_up = "low";

dffeas \delay_signals[2][1] (
	.clk(clk),
	.d(\delay_signals[3][1]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][1]~q ),
	.prn(vcc));
defparam \delay_signals[2][1] .is_wysiwyg = "true";
defparam \delay_signals[2][1] .power_up = "low";

dffeas \delay_signals[1][1] (
	.clk(clk),
	.d(\delay_signals[2][1]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][1]~q ),
	.prn(vcc));
defparam \delay_signals[1][1] .is_wysiwyg = "true";
defparam \delay_signals[1][1] .power_up = "low";

dffeas \delay_signals[3][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][0]~q ),
	.prn(vcc));
defparam \delay_signals[3][0] .is_wysiwyg = "true";
defparam \delay_signals[3][0] .power_up = "low";

dffeas \delay_signals[2][0] (
	.clk(clk),
	.d(\delay_signals[3][0]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][0]~q ),
	.prn(vcc));
defparam \delay_signals[2][0] .is_wysiwyg = "true";
defparam \delay_signals[2][0] .power_up = "low";

dffeas \delay_signals[1][0] (
	.clk(clk),
	.d(\delay_signals[2][0]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][0]~q ),
	.prn(vcc));
defparam \delay_signals[1][0] .is_wysiwyg = "true";
defparam \delay_signals[1][0] .power_up = "low";

dffeas \delay_signals[3][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][11]~q ),
	.prn(vcc));
defparam \delay_signals[3][11] .is_wysiwyg = "true";
defparam \delay_signals[3][11] .power_up = "low";

dffeas \delay_signals[2][11] (
	.clk(clk),
	.d(\delay_signals[3][11]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][11]~q ),
	.prn(vcc));
defparam \delay_signals[2][11] .is_wysiwyg = "true";
defparam \delay_signals[2][11] .power_up = "low";

dffeas \delay_signals[1][11] (
	.clk(clk),
	.d(\delay_signals[2][11]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][11]~q ),
	.prn(vcc));
defparam \delay_signals[1][11] .is_wysiwyg = "true";
defparam \delay_signals[1][11] .power_up = "low";

dffeas \delay_signals[3][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][10]~q ),
	.prn(vcc));
defparam \delay_signals[3][10] .is_wysiwyg = "true";
defparam \delay_signals[3][10] .power_up = "low";

dffeas \delay_signals[2][10] (
	.clk(clk),
	.d(\delay_signals[3][10]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][10]~q ),
	.prn(vcc));
defparam \delay_signals[2][10] .is_wysiwyg = "true";
defparam \delay_signals[2][10] .power_up = "low";

dffeas \delay_signals[1][10] (
	.clk(clk),
	.d(\delay_signals[2][10]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][10]~q ),
	.prn(vcc));
defparam \delay_signals[1][10] .is_wysiwyg = "true";
defparam \delay_signals[1][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_19 (
	aclr,
	delay_signals_7_0,
	delay_signals_9_0,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_10_0,
	delay_signals_11_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_7_0;
output 	delay_signals_9_0;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_10_0;
output 	delay_signals_11_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \delay_signals[1][7]~q ;
wire \delay_signals[1][9]~q ;
wire \delay_signals[1][6]~q ;
wire \delay_signals[1][8]~q ;
wire \delay_signals[1][5]~q ;
wire \delay_signals[1][4]~q ;
wire \delay_signals[1][3]~q ;
wire \delay_signals[1][2]~q ;
wire \delay_signals[1][1]~q ;
wire \delay_signals[1][0]~q ;
wire \delay_signals[1][10]~q ;
wire \delay_signals[1][11]~q ;


dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(\delay_signals[1][7]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(\delay_signals[1][9]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(\delay_signals[1][6]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(\delay_signals[1][8]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(\delay_signals[1][5]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(\delay_signals[1][4]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(\delay_signals[1][3]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(\delay_signals[1][2]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(\delay_signals[1][1]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(\delay_signals[1][0]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(\delay_signals[1][10]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(\delay_signals[1][11]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[1][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][7]~q ),
	.prn(vcc));
defparam \delay_signals[1][7] .is_wysiwyg = "true";
defparam \delay_signals[1][7] .power_up = "low";

dffeas \delay_signals[1][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][9]~q ),
	.prn(vcc));
defparam \delay_signals[1][9] .is_wysiwyg = "true";
defparam \delay_signals[1][9] .power_up = "low";

dffeas \delay_signals[1][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][6]~q ),
	.prn(vcc));
defparam \delay_signals[1][6] .is_wysiwyg = "true";
defparam \delay_signals[1][6] .power_up = "low";

dffeas \delay_signals[1][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][8]~q ),
	.prn(vcc));
defparam \delay_signals[1][8] .is_wysiwyg = "true";
defparam \delay_signals[1][8] .power_up = "low";

dffeas \delay_signals[1][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][5]~q ),
	.prn(vcc));
defparam \delay_signals[1][5] .is_wysiwyg = "true";
defparam \delay_signals[1][5] .power_up = "low";

dffeas \delay_signals[1][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][4]~q ),
	.prn(vcc));
defparam \delay_signals[1][4] .is_wysiwyg = "true";
defparam \delay_signals[1][4] .power_up = "low";

dffeas \delay_signals[1][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][3]~q ),
	.prn(vcc));
defparam \delay_signals[1][3] .is_wysiwyg = "true";
defparam \delay_signals[1][3] .power_up = "low";

dffeas \delay_signals[1][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][2]~q ),
	.prn(vcc));
defparam \delay_signals[1][2] .is_wysiwyg = "true";
defparam \delay_signals[1][2] .power_up = "low";

dffeas \delay_signals[1][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][1]~q ),
	.prn(vcc));
defparam \delay_signals[1][1] .is_wysiwyg = "true";
defparam \delay_signals[1][1] .power_up = "low";

dffeas \delay_signals[1][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][0]~q ),
	.prn(vcc));
defparam \delay_signals[1][0] .is_wysiwyg = "true";
defparam \delay_signals[1][0] .power_up = "low";

dffeas \delay_signals[1][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][10]~q ),
	.prn(vcc));
defparam \delay_signals[1][10] .is_wysiwyg = "true";
defparam \delay_signals[1][10] .power_up = "low";

dffeas \delay_signals[1][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][11]~q ),
	.prn(vcc));
defparam \delay_signals[1][11] .is_wysiwyg = "true";
defparam \delay_signals[1][11] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_20 (
	aclr,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_21 (
	aclr,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	delay_signals_8_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_22 (
	aclr,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_9_0,
	delay_signals_7_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_11_0,
	delay_signals_10_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_9_0;
output 	delay_signals_7_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_23 (
	aclr,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_24 (
	aclr,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_25 (
	aclr,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_26 (
	aclr,
	delay_signals_2_0,
	delay_signals_9_0,
	delay_signals_1_0,
	delay_signals_8_0,
	delay_signals_0_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_10_0,
	delay_signals_11_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_2_0;
output 	delay_signals_9_0;
output 	delay_signals_1_0;
output 	delay_signals_8_0;
output 	delay_signals_0_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_10_0;
output 	delay_signals_11_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_27 (
	aclr,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_28 (
	aclr,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_29 (
	aclr,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_30 (
	aclr,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	delay_signals_8_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_31 (
	aclr,
	u1_m0_wo0_mtree_mult1_8_sub_1_o_1,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	xin,
	delay_signals_11_0,
	delay_signals_10_0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	u1_m0_wo0_mtree_mult1_8_sub_1_o_1;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
input 	[11:0] xin;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \delay_signals[1][9]~q ;
wire \delay_signals[1][8]~q ;
wire \delay_signals[1][7]~q ;
wire \delay_signals[1][6]~q ;
wire \delay_signals[1][5]~q ;
wire \delay_signals[1][4]~q ;
wire \delay_signals[1][3]~q ;
wire \delay_signals[1][2]~q ;
wire \delay_signals[1][11]~q ;
wire \delay_signals[1][10]~q ;


dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(\delay_signals[1][9]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(\delay_signals[1][8]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(\delay_signals[1][7]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(\delay_signals[1][6]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(\delay_signals[1][5]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(\delay_signals[1][4]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(\delay_signals[1][3]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(\delay_signals[1][2]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(u1_m0_wo0_mtree_mult1_8_sub_1_o_1),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(\delay_signals[1][11]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(\delay_signals[1][10]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[1][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][9]~q ),
	.prn(vcc));
defparam \delay_signals[1][9] .is_wysiwyg = "true";
defparam \delay_signals[1][9] .power_up = "low";

dffeas \delay_signals[1][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][8]~q ),
	.prn(vcc));
defparam \delay_signals[1][8] .is_wysiwyg = "true";
defparam \delay_signals[1][8] .power_up = "low";

dffeas \delay_signals[1][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][7]~q ),
	.prn(vcc));
defparam \delay_signals[1][7] .is_wysiwyg = "true";
defparam \delay_signals[1][7] .power_up = "low";

dffeas \delay_signals[1][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][6]~q ),
	.prn(vcc));
defparam \delay_signals[1][6] .is_wysiwyg = "true";
defparam \delay_signals[1][6] .power_up = "low";

dffeas \delay_signals[1][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][5]~q ),
	.prn(vcc));
defparam \delay_signals[1][5] .is_wysiwyg = "true";
defparam \delay_signals[1][5] .power_up = "low";

dffeas \delay_signals[1][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][4]~q ),
	.prn(vcc));
defparam \delay_signals[1][4] .is_wysiwyg = "true";
defparam \delay_signals[1][4] .power_up = "low";

dffeas \delay_signals[1][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][3]~q ),
	.prn(vcc));
defparam \delay_signals[1][3] .is_wysiwyg = "true";
defparam \delay_signals[1][3] .power_up = "low";

dffeas \delay_signals[1][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][2]~q ),
	.prn(vcc));
defparam \delay_signals[1][2] .is_wysiwyg = "true";
defparam \delay_signals[1][2] .power_up = "low";

dffeas \delay_signals[1][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][11]~q ),
	.prn(vcc));
defparam \delay_signals[1][11] .is_wysiwyg = "true";
defparam \delay_signals[1][11] .power_up = "low";

dffeas \delay_signals[1][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][10]~q ),
	.prn(vcc));
defparam \delay_signals[1][10] .is_wysiwyg = "true";
defparam \delay_signals[1][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_32 (
	aclr,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_11_0,
	delay_signals_10_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_33 (
	aclr,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \delay_signals[2][9]~q ;
wire \delay_signals[1][9]~q ;
wire \delay_signals[2][8]~q ;
wire \delay_signals[1][8]~q ;
wire \delay_signals[2][7]~q ;
wire \delay_signals[1][7]~q ;
wire \delay_signals[2][6]~q ;
wire \delay_signals[1][6]~q ;
wire \delay_signals[2][5]~q ;
wire \delay_signals[1][5]~q ;
wire \delay_signals[2][4]~q ;
wire \delay_signals[1][4]~q ;
wire \delay_signals[2][3]~q ;
wire \delay_signals[1][3]~q ;
wire \delay_signals[2][2]~q ;
wire \delay_signals[1][2]~q ;
wire \delay_signals[2][0]~q ;
wire \delay_signals[1][0]~q ;
wire \delay_signals[2][1]~q ;
wire \delay_signals[1][1]~q ;
wire \delay_signals[2][11]~q ;
wire \delay_signals[1][11]~q ;
wire \delay_signals[2][10]~q ;
wire \delay_signals[1][10]~q ;


dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(\delay_signals[1][9]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(\delay_signals[1][8]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(\delay_signals[1][7]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(\delay_signals[1][6]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(\delay_signals[1][5]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(\delay_signals[1][4]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(\delay_signals[1][3]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(\delay_signals[1][2]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(\delay_signals[1][0]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(\delay_signals[1][1]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(\delay_signals[1][11]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(\delay_signals[1][10]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[2][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][9]~q ),
	.prn(vcc));
defparam \delay_signals[2][9] .is_wysiwyg = "true";
defparam \delay_signals[2][9] .power_up = "low";

dffeas \delay_signals[1][9] (
	.clk(clk),
	.d(\delay_signals[2][9]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][9]~q ),
	.prn(vcc));
defparam \delay_signals[1][9] .is_wysiwyg = "true";
defparam \delay_signals[1][9] .power_up = "low";

dffeas \delay_signals[2][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][8]~q ),
	.prn(vcc));
defparam \delay_signals[2][8] .is_wysiwyg = "true";
defparam \delay_signals[2][8] .power_up = "low";

dffeas \delay_signals[1][8] (
	.clk(clk),
	.d(\delay_signals[2][8]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][8]~q ),
	.prn(vcc));
defparam \delay_signals[1][8] .is_wysiwyg = "true";
defparam \delay_signals[1][8] .power_up = "low";

dffeas \delay_signals[2][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][7]~q ),
	.prn(vcc));
defparam \delay_signals[2][7] .is_wysiwyg = "true";
defparam \delay_signals[2][7] .power_up = "low";

dffeas \delay_signals[1][7] (
	.clk(clk),
	.d(\delay_signals[2][7]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][7]~q ),
	.prn(vcc));
defparam \delay_signals[1][7] .is_wysiwyg = "true";
defparam \delay_signals[1][7] .power_up = "low";

dffeas \delay_signals[2][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][6]~q ),
	.prn(vcc));
defparam \delay_signals[2][6] .is_wysiwyg = "true";
defparam \delay_signals[2][6] .power_up = "low";

dffeas \delay_signals[1][6] (
	.clk(clk),
	.d(\delay_signals[2][6]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][6]~q ),
	.prn(vcc));
defparam \delay_signals[1][6] .is_wysiwyg = "true";
defparam \delay_signals[1][6] .power_up = "low";

dffeas \delay_signals[2][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][5]~q ),
	.prn(vcc));
defparam \delay_signals[2][5] .is_wysiwyg = "true";
defparam \delay_signals[2][5] .power_up = "low";

dffeas \delay_signals[1][5] (
	.clk(clk),
	.d(\delay_signals[2][5]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][5]~q ),
	.prn(vcc));
defparam \delay_signals[1][5] .is_wysiwyg = "true";
defparam \delay_signals[1][5] .power_up = "low";

dffeas \delay_signals[2][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][4]~q ),
	.prn(vcc));
defparam \delay_signals[2][4] .is_wysiwyg = "true";
defparam \delay_signals[2][4] .power_up = "low";

dffeas \delay_signals[1][4] (
	.clk(clk),
	.d(\delay_signals[2][4]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][4]~q ),
	.prn(vcc));
defparam \delay_signals[1][4] .is_wysiwyg = "true";
defparam \delay_signals[1][4] .power_up = "low";

dffeas \delay_signals[2][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][3]~q ),
	.prn(vcc));
defparam \delay_signals[2][3] .is_wysiwyg = "true";
defparam \delay_signals[2][3] .power_up = "low";

dffeas \delay_signals[1][3] (
	.clk(clk),
	.d(\delay_signals[2][3]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][3]~q ),
	.prn(vcc));
defparam \delay_signals[1][3] .is_wysiwyg = "true";
defparam \delay_signals[1][3] .power_up = "low";

dffeas \delay_signals[2][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][2]~q ),
	.prn(vcc));
defparam \delay_signals[2][2] .is_wysiwyg = "true";
defparam \delay_signals[2][2] .power_up = "low";

dffeas \delay_signals[1][2] (
	.clk(clk),
	.d(\delay_signals[2][2]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][2]~q ),
	.prn(vcc));
defparam \delay_signals[1][2] .is_wysiwyg = "true";
defparam \delay_signals[1][2] .power_up = "low";

dffeas \delay_signals[2][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][0]~q ),
	.prn(vcc));
defparam \delay_signals[2][0] .is_wysiwyg = "true";
defparam \delay_signals[2][0] .power_up = "low";

dffeas \delay_signals[1][0] (
	.clk(clk),
	.d(\delay_signals[2][0]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][0]~q ),
	.prn(vcc));
defparam \delay_signals[1][0] .is_wysiwyg = "true";
defparam \delay_signals[1][0] .power_up = "low";

dffeas \delay_signals[2][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][1]~q ),
	.prn(vcc));
defparam \delay_signals[2][1] .is_wysiwyg = "true";
defparam \delay_signals[2][1] .power_up = "low";

dffeas \delay_signals[1][1] (
	.clk(clk),
	.d(\delay_signals[2][1]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][1]~q ),
	.prn(vcc));
defparam \delay_signals[1][1] .is_wysiwyg = "true";
defparam \delay_signals[1][1] .power_up = "low";

dffeas \delay_signals[2][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][11]~q ),
	.prn(vcc));
defparam \delay_signals[2][11] .is_wysiwyg = "true";
defparam \delay_signals[2][11] .power_up = "low";

dffeas \delay_signals[1][11] (
	.clk(clk),
	.d(\delay_signals[2][11]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][11]~q ),
	.prn(vcc));
defparam \delay_signals[1][11] .is_wysiwyg = "true";
defparam \delay_signals[1][11] .power_up = "low";

dffeas \delay_signals[2][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][10]~q ),
	.prn(vcc));
defparam \delay_signals[2][10] .is_wysiwyg = "true";
defparam \delay_signals[2][10] .power_up = "low";

dffeas \delay_signals[1][10] (
	.clk(clk),
	.d(\delay_signals[2][10]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][10]~q ),
	.prn(vcc));
defparam \delay_signals[1][10] .is_wysiwyg = "true";
defparam \delay_signals[1][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_34 (
	aclr,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_11_0,
	delay_signals_10_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \delay_signals[3][9]~q ;
wire \delay_signals[2][9]~q ;
wire \delay_signals[1][9]~q ;
wire \delay_signals[3][8]~q ;
wire \delay_signals[2][8]~q ;
wire \delay_signals[1][8]~q ;
wire \delay_signals[3][7]~q ;
wire \delay_signals[2][7]~q ;
wire \delay_signals[1][7]~q ;
wire \delay_signals[3][6]~q ;
wire \delay_signals[2][6]~q ;
wire \delay_signals[1][6]~q ;
wire \delay_signals[3][5]~q ;
wire \delay_signals[2][5]~q ;
wire \delay_signals[1][5]~q ;
wire \delay_signals[3][4]~q ;
wire \delay_signals[2][4]~q ;
wire \delay_signals[1][4]~q ;
wire \delay_signals[3][3]~q ;
wire \delay_signals[2][3]~q ;
wire \delay_signals[1][3]~q ;
wire \delay_signals[3][2]~q ;
wire \delay_signals[2][2]~q ;
wire \delay_signals[1][2]~q ;
wire \delay_signals[3][1]~q ;
wire \delay_signals[2][1]~q ;
wire \delay_signals[1][1]~q ;
wire \delay_signals[3][0]~q ;
wire \delay_signals[2][0]~q ;
wire \delay_signals[1][0]~q ;
wire \delay_signals[3][11]~q ;
wire \delay_signals[2][11]~q ;
wire \delay_signals[1][11]~q ;
wire \delay_signals[3][10]~q ;
wire \delay_signals[2][10]~q ;
wire \delay_signals[1][10]~q ;


dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(\delay_signals[1][9]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(\delay_signals[1][8]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(\delay_signals[1][7]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(\delay_signals[1][6]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(\delay_signals[1][5]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(\delay_signals[1][4]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(\delay_signals[1][3]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(\delay_signals[1][2]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(\delay_signals[1][1]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(\delay_signals[1][0]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(\delay_signals[1][11]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(\delay_signals[1][10]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[3][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][9]~q ),
	.prn(vcc));
defparam \delay_signals[3][9] .is_wysiwyg = "true";
defparam \delay_signals[3][9] .power_up = "low";

dffeas \delay_signals[2][9] (
	.clk(clk),
	.d(\delay_signals[3][9]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][9]~q ),
	.prn(vcc));
defparam \delay_signals[2][9] .is_wysiwyg = "true";
defparam \delay_signals[2][9] .power_up = "low";

dffeas \delay_signals[1][9] (
	.clk(clk),
	.d(\delay_signals[2][9]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][9]~q ),
	.prn(vcc));
defparam \delay_signals[1][9] .is_wysiwyg = "true";
defparam \delay_signals[1][9] .power_up = "low";

dffeas \delay_signals[3][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][8]~q ),
	.prn(vcc));
defparam \delay_signals[3][8] .is_wysiwyg = "true";
defparam \delay_signals[3][8] .power_up = "low";

dffeas \delay_signals[2][8] (
	.clk(clk),
	.d(\delay_signals[3][8]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][8]~q ),
	.prn(vcc));
defparam \delay_signals[2][8] .is_wysiwyg = "true";
defparam \delay_signals[2][8] .power_up = "low";

dffeas \delay_signals[1][8] (
	.clk(clk),
	.d(\delay_signals[2][8]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][8]~q ),
	.prn(vcc));
defparam \delay_signals[1][8] .is_wysiwyg = "true";
defparam \delay_signals[1][8] .power_up = "low";

dffeas \delay_signals[3][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][7]~q ),
	.prn(vcc));
defparam \delay_signals[3][7] .is_wysiwyg = "true";
defparam \delay_signals[3][7] .power_up = "low";

dffeas \delay_signals[2][7] (
	.clk(clk),
	.d(\delay_signals[3][7]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][7]~q ),
	.prn(vcc));
defparam \delay_signals[2][7] .is_wysiwyg = "true";
defparam \delay_signals[2][7] .power_up = "low";

dffeas \delay_signals[1][7] (
	.clk(clk),
	.d(\delay_signals[2][7]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][7]~q ),
	.prn(vcc));
defparam \delay_signals[1][7] .is_wysiwyg = "true";
defparam \delay_signals[1][7] .power_up = "low";

dffeas \delay_signals[3][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][6]~q ),
	.prn(vcc));
defparam \delay_signals[3][6] .is_wysiwyg = "true";
defparam \delay_signals[3][6] .power_up = "low";

dffeas \delay_signals[2][6] (
	.clk(clk),
	.d(\delay_signals[3][6]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][6]~q ),
	.prn(vcc));
defparam \delay_signals[2][6] .is_wysiwyg = "true";
defparam \delay_signals[2][6] .power_up = "low";

dffeas \delay_signals[1][6] (
	.clk(clk),
	.d(\delay_signals[2][6]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][6]~q ),
	.prn(vcc));
defparam \delay_signals[1][6] .is_wysiwyg = "true";
defparam \delay_signals[1][6] .power_up = "low";

dffeas \delay_signals[3][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][5]~q ),
	.prn(vcc));
defparam \delay_signals[3][5] .is_wysiwyg = "true";
defparam \delay_signals[3][5] .power_up = "low";

dffeas \delay_signals[2][5] (
	.clk(clk),
	.d(\delay_signals[3][5]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][5]~q ),
	.prn(vcc));
defparam \delay_signals[2][5] .is_wysiwyg = "true";
defparam \delay_signals[2][5] .power_up = "low";

dffeas \delay_signals[1][5] (
	.clk(clk),
	.d(\delay_signals[2][5]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][5]~q ),
	.prn(vcc));
defparam \delay_signals[1][5] .is_wysiwyg = "true";
defparam \delay_signals[1][5] .power_up = "low";

dffeas \delay_signals[3][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][4]~q ),
	.prn(vcc));
defparam \delay_signals[3][4] .is_wysiwyg = "true";
defparam \delay_signals[3][4] .power_up = "low";

dffeas \delay_signals[2][4] (
	.clk(clk),
	.d(\delay_signals[3][4]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][4]~q ),
	.prn(vcc));
defparam \delay_signals[2][4] .is_wysiwyg = "true";
defparam \delay_signals[2][4] .power_up = "low";

dffeas \delay_signals[1][4] (
	.clk(clk),
	.d(\delay_signals[2][4]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][4]~q ),
	.prn(vcc));
defparam \delay_signals[1][4] .is_wysiwyg = "true";
defparam \delay_signals[1][4] .power_up = "low";

dffeas \delay_signals[3][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][3]~q ),
	.prn(vcc));
defparam \delay_signals[3][3] .is_wysiwyg = "true";
defparam \delay_signals[3][3] .power_up = "low";

dffeas \delay_signals[2][3] (
	.clk(clk),
	.d(\delay_signals[3][3]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][3]~q ),
	.prn(vcc));
defparam \delay_signals[2][3] .is_wysiwyg = "true";
defparam \delay_signals[2][3] .power_up = "low";

dffeas \delay_signals[1][3] (
	.clk(clk),
	.d(\delay_signals[2][3]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][3]~q ),
	.prn(vcc));
defparam \delay_signals[1][3] .is_wysiwyg = "true";
defparam \delay_signals[1][3] .power_up = "low";

dffeas \delay_signals[3][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][2]~q ),
	.prn(vcc));
defparam \delay_signals[3][2] .is_wysiwyg = "true";
defparam \delay_signals[3][2] .power_up = "low";

dffeas \delay_signals[2][2] (
	.clk(clk),
	.d(\delay_signals[3][2]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][2]~q ),
	.prn(vcc));
defparam \delay_signals[2][2] .is_wysiwyg = "true";
defparam \delay_signals[2][2] .power_up = "low";

dffeas \delay_signals[1][2] (
	.clk(clk),
	.d(\delay_signals[2][2]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][2]~q ),
	.prn(vcc));
defparam \delay_signals[1][2] .is_wysiwyg = "true";
defparam \delay_signals[1][2] .power_up = "low";

dffeas \delay_signals[3][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][1]~q ),
	.prn(vcc));
defparam \delay_signals[3][1] .is_wysiwyg = "true";
defparam \delay_signals[3][1] .power_up = "low";

dffeas \delay_signals[2][1] (
	.clk(clk),
	.d(\delay_signals[3][1]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][1]~q ),
	.prn(vcc));
defparam \delay_signals[2][1] .is_wysiwyg = "true";
defparam \delay_signals[2][1] .power_up = "low";

dffeas \delay_signals[1][1] (
	.clk(clk),
	.d(\delay_signals[2][1]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][1]~q ),
	.prn(vcc));
defparam \delay_signals[1][1] .is_wysiwyg = "true";
defparam \delay_signals[1][1] .power_up = "low";

dffeas \delay_signals[3][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][0]~q ),
	.prn(vcc));
defparam \delay_signals[3][0] .is_wysiwyg = "true";
defparam \delay_signals[3][0] .power_up = "low";

dffeas \delay_signals[2][0] (
	.clk(clk),
	.d(\delay_signals[3][0]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][0]~q ),
	.prn(vcc));
defparam \delay_signals[2][0] .is_wysiwyg = "true";
defparam \delay_signals[2][0] .power_up = "low";

dffeas \delay_signals[1][0] (
	.clk(clk),
	.d(\delay_signals[2][0]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][0]~q ),
	.prn(vcc));
defparam \delay_signals[1][0] .is_wysiwyg = "true";
defparam \delay_signals[1][0] .power_up = "low";

dffeas \delay_signals[3][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][11]~q ),
	.prn(vcc));
defparam \delay_signals[3][11] .is_wysiwyg = "true";
defparam \delay_signals[3][11] .power_up = "low";

dffeas \delay_signals[2][11] (
	.clk(clk),
	.d(\delay_signals[3][11]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][11]~q ),
	.prn(vcc));
defparam \delay_signals[2][11] .is_wysiwyg = "true";
defparam \delay_signals[2][11] .power_up = "low";

dffeas \delay_signals[1][11] (
	.clk(clk),
	.d(\delay_signals[2][11]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][11]~q ),
	.prn(vcc));
defparam \delay_signals[1][11] .is_wysiwyg = "true";
defparam \delay_signals[1][11] .power_up = "low";

dffeas \delay_signals[3][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[3][10]~q ),
	.prn(vcc));
defparam \delay_signals[3][10] .is_wysiwyg = "true";
defparam \delay_signals[3][10] .power_up = "low";

dffeas \delay_signals[2][10] (
	.clk(clk),
	.d(\delay_signals[3][10]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[2][10]~q ),
	.prn(vcc));
defparam \delay_signals[2][10] .is_wysiwyg = "true";
defparam \delay_signals[2][10] .power_up = "low";

dffeas \delay_signals[1][10] (
	.clk(clk),
	.d(\delay_signals[2][10]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][10]~q ),
	.prn(vcc));
defparam \delay_signals[1][10] .is_wysiwyg = "true";
defparam \delay_signals[1][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_35 (
	aclr,
	delay_signals_7_0,
	delay_signals_9_0,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_10_0,
	delay_signals_11_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_7_0;
output 	delay_signals_9_0;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_10_0;
output 	delay_signals_11_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \delay_signals[1][7]~q ;
wire \delay_signals[1][9]~q ;
wire \delay_signals[1][6]~q ;
wire \delay_signals[1][8]~q ;
wire \delay_signals[1][5]~q ;
wire \delay_signals[1][4]~q ;
wire \delay_signals[1][3]~q ;
wire \delay_signals[1][2]~q ;
wire \delay_signals[1][1]~q ;
wire \delay_signals[1][0]~q ;
wire \delay_signals[1][10]~q ;
wire \delay_signals[1][11]~q ;


dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(\delay_signals[1][7]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(\delay_signals[1][9]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(\delay_signals[1][6]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(\delay_signals[1][8]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(\delay_signals[1][5]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(\delay_signals[1][4]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(\delay_signals[1][3]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(\delay_signals[1][2]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(\delay_signals[1][1]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(\delay_signals[1][0]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(\delay_signals[1][10]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(\delay_signals[1][11]~q ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[1][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][7]~q ),
	.prn(vcc));
defparam \delay_signals[1][7] .is_wysiwyg = "true";
defparam \delay_signals[1][7] .power_up = "low";

dffeas \delay_signals[1][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][9]~q ),
	.prn(vcc));
defparam \delay_signals[1][9] .is_wysiwyg = "true";
defparam \delay_signals[1][9] .power_up = "low";

dffeas \delay_signals[1][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][6]~q ),
	.prn(vcc));
defparam \delay_signals[1][6] .is_wysiwyg = "true";
defparam \delay_signals[1][6] .power_up = "low";

dffeas \delay_signals[1][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][8]~q ),
	.prn(vcc));
defparam \delay_signals[1][8] .is_wysiwyg = "true";
defparam \delay_signals[1][8] .power_up = "low";

dffeas \delay_signals[1][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][5]~q ),
	.prn(vcc));
defparam \delay_signals[1][5] .is_wysiwyg = "true";
defparam \delay_signals[1][5] .power_up = "low";

dffeas \delay_signals[1][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][4]~q ),
	.prn(vcc));
defparam \delay_signals[1][4] .is_wysiwyg = "true";
defparam \delay_signals[1][4] .power_up = "low";

dffeas \delay_signals[1][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][3]~q ),
	.prn(vcc));
defparam \delay_signals[1][3] .is_wysiwyg = "true";
defparam \delay_signals[1][3] .power_up = "low";

dffeas \delay_signals[1][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][2]~q ),
	.prn(vcc));
defparam \delay_signals[1][2] .is_wysiwyg = "true";
defparam \delay_signals[1][2] .power_up = "low";

dffeas \delay_signals[1][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][1]~q ),
	.prn(vcc));
defparam \delay_signals[1][1] .is_wysiwyg = "true";
defparam \delay_signals[1][1] .power_up = "low";

dffeas \delay_signals[1][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][0]~q ),
	.prn(vcc));
defparam \delay_signals[1][0] .is_wysiwyg = "true";
defparam \delay_signals[1][0] .power_up = "low";

dffeas \delay_signals[1][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][10]~q ),
	.prn(vcc));
defparam \delay_signals[1][10] .is_wysiwyg = "true";
defparam \delay_signals[1][10] .power_up = "low";

dffeas \delay_signals[1][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_signals[1][11]~q ),
	.prn(vcc));
defparam \delay_signals[1][11] .is_wysiwyg = "true";
defparam \delay_signals[1][11] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_36 (
	aclr,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_37 (
	aclr,
	ena,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	ena;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_38 (
	aclr,
	delay_signals_7_0,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	xin,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_7_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
input 	[11:0] xin;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_39 (
	aclr,
	xin,
	ena,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_9_0,
	delay_signals_7_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_11_0,
	delay_signals_10_0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	[11:0] xin;
input 	ena;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_9_0;
output 	delay_signals_7_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_40 (
	aclr,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_9_0,
	delay_signals_7_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_9_0;
output 	delay_signals_7_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_41 (
	aclr,
	delay_signals_4_0,
	delay_signals_6_0,
	delay_signals_9_0,
	delay_signals_5_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	xin,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_4_0;
output 	delay_signals_6_0;
output 	delay_signals_9_0;
output 	delay_signals_5_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
input 	[11:0] xin;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_42 (
	aclr,
	delay_signals_4_0,
	delay_signals_7_0,
	delay_signals_9_0,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_5_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	xin,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_4_0;
output 	delay_signals_7_0;
output 	delay_signals_9_0;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_5_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
input 	[11:0] xin;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_43 (
	aclr,
	delay_signals_2_0,
	delay_signals_9_0,
	delay_signals_1_0,
	delay_signals_8_0,
	delay_signals_0_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	xin,
	delay_signals_10_0,
	delay_signals_11_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_2_0;
output 	delay_signals_9_0;
output 	delay_signals_1_0;
output 	delay_signals_8_0;
output 	delay_signals_0_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
input 	[11:0] xin;
output 	delay_signals_10_0;
output 	delay_signals_11_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_44 (
	aclr,
	delay_signals_4_0,
	delay_signals_7_0,
	delay_signals_9_0,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_5_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	xin,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_4_0;
output 	delay_signals_7_0;
output 	delay_signals_9_0;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_5_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
input 	[11:0] xin;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_45 (
	aclr,
	delay_signals_4_0,
	delay_signals_6_0,
	delay_signals_9_0,
	delay_signals_5_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	xin,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_4_0;
output 	delay_signals_6_0;
output 	delay_signals_9_0;
output 	delay_signals_5_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
input 	[11:0] xin;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_46 (
	aclr,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_9_0,
	delay_signals_7_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	xin,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_9_0;
output 	delay_signals_7_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
input 	[11:0] xin;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_47 (
	aclr,
	xin,
	ena,
	delay_signals_7_0,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	[11:0] xin;
input 	ena;
output 	delay_signals_7_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_48 (
	aclr,
	ena,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	ena;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_49 (
	aclr,
	delay_signals_7_0,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_7_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_50 (
	aclr,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	xin,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
input 	[11:0] xin;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_51 (
	aclr,
	delay_signals_7_0,
	delay_signals_9_0,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	xin,
	delay_signals_10_0,
	delay_signals_11_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_7_0;
output 	delay_signals_9_0;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
input 	[11:0] xin;
output 	delay_signals_10_0;
output 	delay_signals_11_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_52 (
	aclr,
	xin,
	ena,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_11_0,
	delay_signals_10_0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	[11:0] xin;
input 	ena;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_53 (
	aclr,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_54 (
	aclr,
	xin,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	[11:0] xin;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_55 (
	aclr,
	ena,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	ena;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_56 (
	aclr,
	ena,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	ena;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_57 (
	aclr,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_58 (
	aclr,
	delay_signals_9_0,
	xin,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_9_0;
input 	[11:0] xin;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_59 (
	aclr,
	xin,
	ena,
	delay_signals_7_0,
	delay_signals_9_0,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_10_0,
	delay_signals_11_0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	[11:0] xin;
input 	ena;
output 	delay_signals_7_0;
output 	delay_signals_9_0;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_10_0;
output 	delay_signals_11_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_60 (
	aclr,
	delay_signals_7_0,
	delay_signals_9_0,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_10_0,
	delay_signals_11_0,
	ena,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_7_0;
output 	delay_signals_9_0;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_10_0;
output 	delay_signals_11_0;
input 	ena;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_61 (
	aclr,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	xin,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
input 	[11:0] xin;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_62 (
	aclr,
	ena,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	ena;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_63 (
	aclr,
	delay_signals_7_0,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	xin,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_7_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
input 	[11:0] xin;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_64 (
	aclr,
	xin,
	ena,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_9_0,
	delay_signals_7_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_11_0,
	delay_signals_10_0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	[11:0] xin;
input 	ena;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_9_0;
output 	delay_signals_7_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_65 (
	aclr,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_9_0,
	delay_signals_7_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_9_0;
output 	delay_signals_7_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_66 (
	aclr,
	delay_signals_4_0,
	delay_signals_6_0,
	delay_signals_9_0,
	delay_signals_5_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	xin,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_4_0;
output 	delay_signals_6_0;
output 	delay_signals_9_0;
output 	delay_signals_5_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
input 	[11:0] xin;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_67 (
	aclr,
	delay_signals_4_0,
	delay_signals_7_0,
	delay_signals_9_0,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_5_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	xin,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_4_0;
output 	delay_signals_7_0;
output 	delay_signals_9_0;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_5_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
input 	[11:0] xin;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_68 (
	aclr,
	delay_signals_2_0,
	delay_signals_9_0,
	delay_signals_1_0,
	delay_signals_8_0,
	delay_signals_0_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	xin,
	delay_signals_10_0,
	delay_signals_11_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_2_0;
output 	delay_signals_9_0;
output 	delay_signals_1_0;
output 	delay_signals_8_0;
output 	delay_signals_0_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
input 	[11:0] xin;
output 	delay_signals_10_0;
output 	delay_signals_11_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_69 (
	aclr,
	delay_signals_4_0,
	delay_signals_7_0,
	delay_signals_9_0,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_5_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	xin,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_4_0;
output 	delay_signals_7_0;
output 	delay_signals_9_0;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_5_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
input 	[11:0] xin;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_70 (
	aclr,
	delay_signals_4_0,
	delay_signals_6_0,
	delay_signals_9_0,
	delay_signals_5_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	xin,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_4_0;
output 	delay_signals_6_0;
output 	delay_signals_9_0;
output 	delay_signals_5_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
input 	[11:0] xin;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_71 (
	aclr,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_9_0,
	delay_signals_7_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	xin,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_9_0;
output 	delay_signals_7_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
input 	[11:0] xin;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_72 (
	aclr,
	xin,
	ena,
	delay_signals_7_0,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	[11:0] xin;
input 	ena;
output 	delay_signals_7_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_73 (
	aclr,
	ena,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	ena;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_74 (
	aclr,
	delay_signals_7_0,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_7_0;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_75 (
	aclr,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	xin,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
input 	[11:0] xin;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_76 (
	aclr,
	delay_signals_7_0,
	delay_signals_9_0,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	xin,
	delay_signals_10_0,
	delay_signals_11_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_7_0;
output 	delay_signals_9_0;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
input 	[11:0] xin;
output 	delay_signals_10_0;
output 	delay_signals_11_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_77 (
	aclr,
	xin,
	ena,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_11_0,
	delay_signals_10_0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	[11:0] xin;
input 	ena;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_78 (
	aclr,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_79 (
	aclr,
	xin,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	[11:0] xin;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_80 (
	aclr,
	ena,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	ena;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_81 (
	aclr,
	ena,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	ena;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_82 (
	aclr,
	delay_signals_9_0,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_0_0,
	delay_signals_1_0,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_9_0;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_0_0;
output 	delay_signals_1_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_83 (
	aclr,
	delay_signals_9_0,
	xin,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_11_0,
	delay_signals_10_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_9_0;
input 	[11:0] xin;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_84 (
	aclr,
	xin,
	ena,
	delay_signals_7_0,
	delay_signals_9_0,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_10_0,
	delay_signals_11_0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
input 	[11:0] xin;
input 	ena;
output 	delay_signals_7_0;
output 	delay_signals_9_0;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_10_0;
output 	delay_signals_11_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_85 (
	aclr,
	delay_signals_7_0,
	delay_signals_9_0,
	delay_signals_6_0,
	delay_signals_8_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	delay_signals_10_0,
	delay_signals_11_0,
	ena,
	xin,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_7_0;
output 	delay_signals_9_0;
output 	delay_signals_6_0;
output 	delay_signals_8_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
output 	delay_signals_10_0;
output 	delay_signals_11_0;
input 	ena;
input 	[11:0] xin;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

endmodule

module lms_dsp_dspba_delay_86 (
	aclr,
	delay_signals_8_0,
	delay_signals_7_0,
	delay_signals_6_0,
	delay_signals_5_0,
	delay_signals_4_0,
	delay_signals_3_0,
	delay_signals_2_0,
	delay_signals_1_0,
	delay_signals_0_0,
	xin,
	delay_signals_11_0,
	delay_signals_10_0,
	delay_signals_9_0,
	ena,
	clk)/* synthesis synthesis_greybox=0 */;
input 	aclr;
output 	delay_signals_8_0;
output 	delay_signals_7_0;
output 	delay_signals_6_0;
output 	delay_signals_5_0;
output 	delay_signals_4_0;
output 	delay_signals_3_0;
output 	delay_signals_2_0;
output 	delay_signals_1_0;
output 	delay_signals_0_0;
input 	[11:0] xin;
output 	delay_signals_11_0;
output 	delay_signals_10_0;
output 	delay_signals_9_0;
input 	ena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \delay_signals[0][8] (
	.clk(clk),
	.d(xin[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_8_0),
	.prn(vcc));
defparam \delay_signals[0][8] .is_wysiwyg = "true";
defparam \delay_signals[0][8] .power_up = "low";

dffeas \delay_signals[0][7] (
	.clk(clk),
	.d(xin[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_7_0),
	.prn(vcc));
defparam \delay_signals[0][7] .is_wysiwyg = "true";
defparam \delay_signals[0][7] .power_up = "low";

dffeas \delay_signals[0][6] (
	.clk(clk),
	.d(xin[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_6_0),
	.prn(vcc));
defparam \delay_signals[0][6] .is_wysiwyg = "true";
defparam \delay_signals[0][6] .power_up = "low";

dffeas \delay_signals[0][5] (
	.clk(clk),
	.d(xin[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_5_0),
	.prn(vcc));
defparam \delay_signals[0][5] .is_wysiwyg = "true";
defparam \delay_signals[0][5] .power_up = "low";

dffeas \delay_signals[0][4] (
	.clk(clk),
	.d(xin[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_4_0),
	.prn(vcc));
defparam \delay_signals[0][4] .is_wysiwyg = "true";
defparam \delay_signals[0][4] .power_up = "low";

dffeas \delay_signals[0][3] (
	.clk(clk),
	.d(xin[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_3_0),
	.prn(vcc));
defparam \delay_signals[0][3] .is_wysiwyg = "true";
defparam \delay_signals[0][3] .power_up = "low";

dffeas \delay_signals[0][2] (
	.clk(clk),
	.d(xin[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_2_0),
	.prn(vcc));
defparam \delay_signals[0][2] .is_wysiwyg = "true";
defparam \delay_signals[0][2] .power_up = "low";

dffeas \delay_signals[0][1] (
	.clk(clk),
	.d(xin[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_1_0),
	.prn(vcc));
defparam \delay_signals[0][1] .is_wysiwyg = "true";
defparam \delay_signals[0][1] .power_up = "low";

dffeas \delay_signals[0][0] (
	.clk(clk),
	.d(xin[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_0_0),
	.prn(vcc));
defparam \delay_signals[0][0] .is_wysiwyg = "true";
defparam \delay_signals[0][0] .power_up = "low";

dffeas \delay_signals[0][11] (
	.clk(clk),
	.d(xin[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_11_0),
	.prn(vcc));
defparam \delay_signals[0][11] .is_wysiwyg = "true";
defparam \delay_signals[0][11] .power_up = "low";

dffeas \delay_signals[0][10] (
	.clk(clk),
	.d(xin[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_10_0),
	.prn(vcc));
defparam \delay_signals[0][10] .is_wysiwyg = "true";
defparam \delay_signals[0][10] .power_up = "low";

dffeas \delay_signals[0][9] (
	.clk(clk),
	.d(xin[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena),
	.q(delay_signals_9_0),
	.prn(vcc));
defparam \delay_signals[0][9] .is_wysiwyg = "true";
defparam \delay_signals[0][9] .power_up = "low";

endmodule

module lms_dsp_packet_presence_detection (
	count_reg_0,
	short_sum_reg_0,
	short_sum_reg_1,
	short_sum_reg_2,
	short_sum_reg_3,
	short_sum_reg_4,
	short_sum_reg_5,
	short_sum_reg_6,
	short_sum_reg_7,
	short_sum_reg_8,
	short_sum_reg_9,
	short_sum_reg_10,
	short_sum_reg_11,
	short_sum_reg_12,
	short_sum_reg_13,
	short_sum_reg_14,
	short_sum_reg_15,
	short_sum_reg_16,
	short_sum_reg_17,
	count_reg_1,
	count_reg_2,
	count_reg_3,
	count_reg_4,
	count_reg_5,
	count_reg_6,
	count_reg_7,
	count_reg_8,
	count_reg_9,
	count_reg_10,
	count_reg_11,
	count_reg_12,
	count_reg_13,
	count_reg_14,
	count_reg_15,
	long_shift_rescale_0,
	long_shift_rescale_1,
	long_shift_rescale_2,
	long_shift_rescale_3,
	long_shift_rescale_4,
	long_shift_rescale_5,
	long_shift_rescale_6,
	long_shift_rescale_7,
	long_shift_rescale_8,
	long_shift_rescale_9,
	long_shift_rescale_10,
	long_shift_rescale_11,
	long_shift_rescale_12,
	long_shift_rescale_13,
	long_shift_rescale_14,
	long_shift_rescale_15,
	long_shift_rescale_16,
	long_shift_rescale_17,
	long_shift_rescale_18,
	long_shift_rescale_19,
	long_shift_rescale_20,
	altera_reset_synchronizer_int_chain_out,
	data_out_12,
	data_out_0,
	data_out_11,
	data_out_10,
	data_out_9,
	data_out_8,
	data_out_7,
	data_out_6,
	data_out_5,
	data_out_4,
	data_out_3,
	data_out_2,
	data_out_1,
	data_out_23,
	data_out_22,
	data_out_21,
	data_out_20,
	data_out_19,
	data_out_18,
	data_out_17,
	data_out_16,
	data_out_15,
	data_out_14,
	data_out_13,
	data_valid,
	avalon_streaming_source_data_0,
	avalon_streaming_source_data_1,
	avalon_streaming_source_data_2,
	avalon_streaming_source_data_3,
	avalon_streaming_source_data_4,
	avalon_streaming_source_data_5,
	avalon_streaming_source_data_6,
	avalon_streaming_source_data_7,
	avalon_streaming_source_data_8,
	avalon_streaming_source_data_9,
	avalon_streaming_source_data_10,
	avalon_streaming_source_data_11,
	avalon_streaming_source_data_12,
	avalon_streaming_source_data_13,
	avalon_streaming_source_data_14,
	avalon_streaming_source_data_15,
	avalon_streaming_source_data_16,
	avalon_streaming_source_data_17,
	avalon_streaming_source_data_18,
	avalon_streaming_source_data_19,
	avalon_streaming_source_data_20,
	avalon_streaming_source_data_21,
	avalon_streaming_source_data_22,
	avalon_streaming_source_data_23,
	delay_reg_24_3,
	GND_port,
	clk_clk,
	ppd_cfg_passthrough_len_15,
	ppd_cfg_passthrough_len_14,
	ppd_cfg_passthrough_len_13,
	ppd_cfg_passthrough_len_12,
	ppd_cfg_passthrough_len_11,
	ppd_cfg_passthrough_len_10,
	ppd_cfg_passthrough_len_9,
	ppd_cfg_passthrough_len_8,
	ppd_cfg_passthrough_len_7,
	ppd_cfg_passthrough_len_6,
	ppd_cfg_passthrough_len_5,
	ppd_cfg_passthrough_len_4,
	ppd_cfg_passthrough_len_3,
	ppd_cfg_passthrough_len_2,
	ppd_cfg_passthrough_len_1,
	ppd_cfg_passthrough_len_0,
	ppd_cfg_clear_rs,
	ppd_cfg_threshold_0,
	ppd_cfg_threshold_1,
	ppd_cfg_threshold_2,
	ppd_cfg_threshold_3,
	ppd_cfg_threshold_4,
	ppd_cfg_threshold_5,
	ppd_cfg_threshold_6,
	ppd_cfg_threshold_7,
	ppd_cfg_enable)/* synthesis synthesis_greybox=0 */;
output 	count_reg_0;
output 	short_sum_reg_0;
output 	short_sum_reg_1;
output 	short_sum_reg_2;
output 	short_sum_reg_3;
output 	short_sum_reg_4;
output 	short_sum_reg_5;
output 	short_sum_reg_6;
output 	short_sum_reg_7;
output 	short_sum_reg_8;
output 	short_sum_reg_9;
output 	short_sum_reg_10;
output 	short_sum_reg_11;
output 	short_sum_reg_12;
output 	short_sum_reg_13;
output 	short_sum_reg_14;
output 	short_sum_reg_15;
output 	short_sum_reg_16;
output 	short_sum_reg_17;
output 	count_reg_1;
output 	count_reg_2;
output 	count_reg_3;
output 	count_reg_4;
output 	count_reg_5;
output 	count_reg_6;
output 	count_reg_7;
output 	count_reg_8;
output 	count_reg_9;
output 	count_reg_10;
output 	count_reg_11;
output 	count_reg_12;
output 	count_reg_13;
output 	count_reg_14;
output 	count_reg_15;
output 	long_shift_rescale_0;
output 	long_shift_rescale_1;
output 	long_shift_rescale_2;
output 	long_shift_rescale_3;
output 	long_shift_rescale_4;
output 	long_shift_rescale_5;
output 	long_shift_rescale_6;
output 	long_shift_rescale_7;
output 	long_shift_rescale_8;
output 	long_shift_rescale_9;
output 	long_shift_rescale_10;
output 	long_shift_rescale_11;
output 	long_shift_rescale_12;
output 	long_shift_rescale_13;
output 	long_shift_rescale_14;
output 	long_shift_rescale_15;
output 	long_shift_rescale_16;
output 	long_shift_rescale_17;
output 	long_shift_rescale_18;
output 	long_shift_rescale_19;
output 	long_shift_rescale_20;
input 	altera_reset_synchronizer_int_chain_out;
input 	data_out_12;
input 	data_out_0;
input 	data_out_11;
input 	data_out_10;
input 	data_out_9;
input 	data_out_8;
input 	data_out_7;
input 	data_out_6;
input 	data_out_5;
input 	data_out_4;
input 	data_out_3;
input 	data_out_2;
input 	data_out_1;
input 	data_out_23;
input 	data_out_22;
input 	data_out_21;
input 	data_out_20;
input 	data_out_19;
input 	data_out_18;
input 	data_out_17;
input 	data_out_16;
input 	data_out_15;
input 	data_out_14;
input 	data_out_13;
input 	data_valid;
output 	avalon_streaming_source_data_0;
output 	avalon_streaming_source_data_1;
output 	avalon_streaming_source_data_2;
output 	avalon_streaming_source_data_3;
output 	avalon_streaming_source_data_4;
output 	avalon_streaming_source_data_5;
output 	avalon_streaming_source_data_6;
output 	avalon_streaming_source_data_7;
output 	avalon_streaming_source_data_8;
output 	avalon_streaming_source_data_9;
output 	avalon_streaming_source_data_10;
output 	avalon_streaming_source_data_11;
output 	avalon_streaming_source_data_12;
output 	avalon_streaming_source_data_13;
output 	avalon_streaming_source_data_14;
output 	avalon_streaming_source_data_15;
output 	avalon_streaming_source_data_16;
output 	avalon_streaming_source_data_17;
output 	avalon_streaming_source_data_18;
output 	avalon_streaming_source_data_19;
output 	avalon_streaming_source_data_20;
output 	avalon_streaming_source_data_21;
output 	avalon_streaming_source_data_22;
output 	avalon_streaming_source_data_23;
output 	delay_reg_24_3;
input 	GND_port;
input 	clk_clk;
input 	ppd_cfg_passthrough_len_15;
input 	ppd_cfg_passthrough_len_14;
input 	ppd_cfg_passthrough_len_13;
input 	ppd_cfg_passthrough_len_12;
input 	ppd_cfg_passthrough_len_11;
input 	ppd_cfg_passthrough_len_10;
input 	ppd_cfg_passthrough_len_9;
input 	ppd_cfg_passthrough_len_8;
input 	ppd_cfg_passthrough_len_7;
input 	ppd_cfg_passthrough_len_6;
input 	ppd_cfg_passthrough_len_5;
input 	ppd_cfg_passthrough_len_4;
input 	ppd_cfg_passthrough_len_3;
input 	ppd_cfg_passthrough_len_2;
input 	ppd_cfg_passthrough_len_1;
input 	ppd_cfg_passthrough_len_0;
input 	ppd_cfg_clear_rs;
input 	ppd_cfg_threshold_0;
input 	ppd_cfg_threshold_1;
input 	ppd_cfg_threshold_2;
input 	ppd_cfg_threshold_3;
input 	ppd_cfg_threshold_4;
input 	ppd_cfg_threshold_5;
input 	ppd_cfg_threshold_6;
input 	ppd_cfg_threshold_7;
input 	ppd_cfg_enable;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \running_sum_inst|LessThan0~34_combout ;
wire \cmplx2mag_inst|mag_reg[0]~q ;
wire \counter_inst|running_reg~q ;
wire \cmplx2mag_inst|mag_reg[1]~q ;
wire \cmplx2mag_inst|mag_reg[2]~q ;
wire \cmplx2mag_inst|mag_reg[3]~q ;
wire \cmplx2mag_inst|mag_reg[4]~q ;
wire \cmplx2mag_inst|mag_reg[5]~q ;
wire \cmplx2mag_inst|mag_reg[6]~q ;
wire \cmplx2mag_inst|mag_reg[7]~q ;
wire \cmplx2mag_inst|mag_reg[8]~q ;
wire \cmplx2mag_inst|mag_reg[9]~q ;
wire \cmplx2mag_inst|mag_reg[10]~q ;
wire \cmplx2mag_inst|mag_reg[11]~q ;
wire \cmplx2mag_inst|mag_reg[12]~q ;
wire \running_sum_inst|launch~2_combout ;
wire \running_sum_inst|long_shift_rescale[25]~q ;
wire \running_sum_inst|launch~combout ;
wire \delay_line_inst|delay_reg[1][24]~q ;
wire \delay_line_inst|delay_reg[0][24]~q ;
wire \delay_line_inst|delay_reg[2][25]~q ;
wire \delay_line_inst|delay_reg[3][0]~q ;
wire \delay_line_inst|delay_reg[3][1]~q ;
wire \delay_line_inst|delay_reg[3][2]~q ;
wire \delay_line_inst|delay_reg[3][3]~q ;
wire \delay_line_inst|delay_reg[3][4]~q ;
wire \delay_line_inst|delay_reg[3][5]~q ;
wire \delay_line_inst|delay_reg[3][6]~q ;
wire \delay_line_inst|delay_reg[3][7]~q ;
wire \delay_line_inst|delay_reg[3][8]~q ;
wire \delay_line_inst|delay_reg[3][9]~q ;
wire \delay_line_inst|delay_reg[3][10]~q ;
wire \delay_line_inst|delay_reg[3][11]~q ;
wire \delay_line_inst|delay_reg[3][12]~q ;
wire \delay_line_inst|delay_reg[3][13]~q ;
wire \delay_line_inst|delay_reg[3][14]~q ;
wire \delay_line_inst|delay_reg[3][15]~q ;
wire \delay_line_inst|delay_reg[3][16]~q ;
wire \delay_line_inst|delay_reg[3][17]~q ;
wire \delay_line_inst|delay_reg[3][18]~q ;
wire \delay_line_inst|delay_reg[3][19]~q ;
wire \delay_line_inst|delay_reg[3][20]~q ;
wire \delay_line_inst|delay_reg[3][21]~q ;
wire \delay_line_inst|delay_reg[3][22]~q ;
wire \delay_line_inst|delay_reg[3][23]~q ;
wire \avalon_streaming_source_data~0_combout ;


lms_dsp_counter counter_inst(
	.count_reg_0(count_reg_0),
	.running_reg1(\counter_inst|running_reg~q ),
	.count_reg_1(count_reg_1),
	.count_reg_2(count_reg_2),
	.count_reg_3(count_reg_3),
	.count_reg_4(count_reg_4),
	.count_reg_5(count_reg_5),
	.count_reg_6(count_reg_6),
	.count_reg_7(count_reg_7),
	.count_reg_8(count_reg_8),
	.count_reg_9(count_reg_9),
	.count_reg_10(count_reg_10),
	.count_reg_11(count_reg_11),
	.count_reg_12(count_reg_12),
	.count_reg_13(count_reg_13),
	.count_reg_14(count_reg_14),
	.count_reg_15(count_reg_15),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.launch(\running_sum_inst|launch~combout ),
	.delay_reg_24_1(\delay_line_inst|delay_reg[1][24]~q ),
	.clock(clk_clk),
	.ppd_cfg_passthrough_len_15(ppd_cfg_passthrough_len_15),
	.ppd_cfg_passthrough_len_14(ppd_cfg_passthrough_len_14),
	.ppd_cfg_passthrough_len_13(ppd_cfg_passthrough_len_13),
	.ppd_cfg_passthrough_len_12(ppd_cfg_passthrough_len_12),
	.ppd_cfg_passthrough_len_11(ppd_cfg_passthrough_len_11),
	.ppd_cfg_passthrough_len_10(ppd_cfg_passthrough_len_10),
	.ppd_cfg_passthrough_len_9(ppd_cfg_passthrough_len_9),
	.ppd_cfg_passthrough_len_8(ppd_cfg_passthrough_len_8),
	.ppd_cfg_passthrough_len_7(ppd_cfg_passthrough_len_7),
	.ppd_cfg_passthrough_len_6(ppd_cfg_passthrough_len_6),
	.ppd_cfg_passthrough_len_5(ppd_cfg_passthrough_len_5),
	.ppd_cfg_passthrough_len_4(ppd_cfg_passthrough_len_4),
	.ppd_cfg_passthrough_len_3(ppd_cfg_passthrough_len_3),
	.ppd_cfg_passthrough_len_2(ppd_cfg_passthrough_len_2),
	.ppd_cfg_passthrough_len_1(ppd_cfg_passthrough_len_1),
	.ppd_cfg_passthrough_len_0(ppd_cfg_passthrough_len_0));

lms_dsp_dual_running_sum running_sum_inst(
	.short_sum_reg_0(short_sum_reg_0),
	.short_sum_reg_1(short_sum_reg_1),
	.short_sum_reg_2(short_sum_reg_2),
	.short_sum_reg_3(short_sum_reg_3),
	.short_sum_reg_4(short_sum_reg_4),
	.short_sum_reg_5(short_sum_reg_5),
	.short_sum_reg_6(short_sum_reg_6),
	.short_sum_reg_7(short_sum_reg_7),
	.short_sum_reg_8(short_sum_reg_8),
	.short_sum_reg_9(short_sum_reg_9),
	.short_sum_reg_10(short_sum_reg_10),
	.short_sum_reg_11(short_sum_reg_11),
	.short_sum_reg_12(short_sum_reg_12),
	.short_sum_reg_13(short_sum_reg_13),
	.short_sum_reg_14(short_sum_reg_14),
	.short_sum_reg_15(short_sum_reg_15),
	.short_sum_reg_16(short_sum_reg_16),
	.short_sum_reg_17(short_sum_reg_17),
	.LessThan0(\running_sum_inst|LessThan0~34_combout ),
	.mag_reg_0(\cmplx2mag_inst|mag_reg[0]~q ),
	.running_reg(\counter_inst|running_reg~q ),
	.mag_reg_1(\cmplx2mag_inst|mag_reg[1]~q ),
	.mag_reg_2(\cmplx2mag_inst|mag_reg[2]~q ),
	.mag_reg_3(\cmplx2mag_inst|mag_reg[3]~q ),
	.mag_reg_4(\cmplx2mag_inst|mag_reg[4]~q ),
	.mag_reg_5(\cmplx2mag_inst|mag_reg[5]~q ),
	.mag_reg_6(\cmplx2mag_inst|mag_reg[6]~q ),
	.mag_reg_7(\cmplx2mag_inst|mag_reg[7]~q ),
	.mag_reg_8(\cmplx2mag_inst|mag_reg[8]~q ),
	.mag_reg_9(\cmplx2mag_inst|mag_reg[9]~q ),
	.mag_reg_10(\cmplx2mag_inst|mag_reg[10]~q ),
	.mag_reg_11(\cmplx2mag_inst|mag_reg[11]~q ),
	.mag_reg_12(\cmplx2mag_inst|mag_reg[12]~q ),
	.long_shift_rescale_0(long_shift_rescale_0),
	.long_shift_rescale_1(long_shift_rescale_1),
	.long_shift_rescale_2(long_shift_rescale_2),
	.long_shift_rescale_3(long_shift_rescale_3),
	.long_shift_rescale_4(long_shift_rescale_4),
	.long_shift_rescale_5(long_shift_rescale_5),
	.long_shift_rescale_6(long_shift_rescale_6),
	.long_shift_rescale_7(long_shift_rescale_7),
	.long_shift_rescale_8(long_shift_rescale_8),
	.long_shift_rescale_9(long_shift_rescale_9),
	.long_shift_rescale_10(long_shift_rescale_10),
	.long_shift_rescale_11(long_shift_rescale_11),
	.long_shift_rescale_12(long_shift_rescale_12),
	.long_shift_rescale_13(long_shift_rescale_13),
	.long_shift_rescale_14(long_shift_rescale_14),
	.long_shift_rescale_15(long_shift_rescale_15),
	.long_shift_rescale_16(long_shift_rescale_16),
	.long_shift_rescale_17(long_shift_rescale_17),
	.long_shift_rescale_18(long_shift_rescale_18),
	.long_shift_rescale_19(long_shift_rescale_19),
	.long_shift_rescale_20(long_shift_rescale_20),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.launch1(\running_sum_inst|launch~2_combout ),
	.long_shift_rescale_25(\running_sum_inst|long_shift_rescale[25]~q ),
	.launch2(\running_sum_inst|launch~combout ),
	.delay_reg_24_0(\delay_line_inst|delay_reg[0][24]~q ),
	.GND_port(GND_port),
	.clk_clk(clk_clk),
	.ppd_cfg_clear_rs(ppd_cfg_clear_rs),
	.ppd_cfg_threshold_0(ppd_cfg_threshold_0),
	.ppd_cfg_threshold_1(ppd_cfg_threshold_1),
	.ppd_cfg_threshold_2(ppd_cfg_threshold_2),
	.ppd_cfg_threshold_3(ppd_cfg_threshold_3),
	.ppd_cfg_threshold_4(ppd_cfg_threshold_4),
	.ppd_cfg_threshold_5(ppd_cfg_threshold_5),
	.ppd_cfg_threshold_6(ppd_cfg_threshold_6),
	.ppd_cfg_threshold_7(ppd_cfg_threshold_7));

lms_dsp_cmplx2mag cmplx2mag_inst(
	.mag_reg_0(\cmplx2mag_inst|mag_reg[0]~q ),
	.mag_reg_1(\cmplx2mag_inst|mag_reg[1]~q ),
	.mag_reg_2(\cmplx2mag_inst|mag_reg[2]~q ),
	.mag_reg_3(\cmplx2mag_inst|mag_reg[3]~q ),
	.mag_reg_4(\cmplx2mag_inst|mag_reg[4]~q ),
	.mag_reg_5(\cmplx2mag_inst|mag_reg[5]~q ),
	.mag_reg_6(\cmplx2mag_inst|mag_reg[6]~q ),
	.mag_reg_7(\cmplx2mag_inst|mag_reg[7]~q ),
	.mag_reg_8(\cmplx2mag_inst|mag_reg[8]~q ),
	.mag_reg_9(\cmplx2mag_inst|mag_reg[9]~q ),
	.mag_reg_10(\cmplx2mag_inst|mag_reg[10]~q ),
	.mag_reg_11(\cmplx2mag_inst|mag_reg[11]~q ),
	.mag_reg_12(\cmplx2mag_inst|mag_reg[12]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.data_out_12(data_out_12),
	.data_out_0(data_out_0),
	.data_out_11(data_out_11),
	.data_out_10(data_out_10),
	.data_out_9(data_out_9),
	.data_out_8(data_out_8),
	.data_out_7(data_out_7),
	.data_out_6(data_out_6),
	.data_out_5(data_out_5),
	.data_out_4(data_out_4),
	.data_out_3(data_out_3),
	.data_out_2(data_out_2),
	.data_out_1(data_out_1),
	.data_out_23(data_out_23),
	.data_out_22(data_out_22),
	.data_out_21(data_out_21),
	.data_out_20(data_out_20),
	.data_out_19(data_out_19),
	.data_out_18(data_out_18),
	.data_out_17(data_out_17),
	.data_out_16(data_out_16),
	.data_out_15(data_out_15),
	.data_out_14(data_out_14),
	.data_out_13(data_out_13),
	.clock(clk_clk));

lms_dsp_delay_line delay_line_inst(
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.delay_reg_24_1(\delay_line_inst|delay_reg[1][24]~q ),
	.delay_reg_24_0(\delay_line_inst|delay_reg[0][24]~q ),
	.data_out_12(data_out_12),
	.data_out_0(data_out_0),
	.data_out_11(data_out_11),
	.data_out_10(data_out_10),
	.data_out_9(data_out_9),
	.data_out_8(data_out_8),
	.data_out_7(data_out_7),
	.data_out_6(data_out_6),
	.data_out_5(data_out_5),
	.data_out_4(data_out_4),
	.data_out_3(data_out_3),
	.data_out_2(data_out_2),
	.data_out_1(data_out_1),
	.data_out_23(data_out_23),
	.data_out_22(data_out_22),
	.data_out_21(data_out_21),
	.data_out_20(data_out_20),
	.data_out_19(data_out_19),
	.data_out_18(data_out_18),
	.data_out_17(data_out_17),
	.data_out_16(data_out_16),
	.data_out_15(data_out_15),
	.data_out_14(data_out_14),
	.data_out_13(data_out_13),
	.data_valid(data_valid),
	.delay_reg_25_2(\delay_line_inst|delay_reg[2][25]~q ),
	.delay_reg_0_3(\delay_line_inst|delay_reg[3][0]~q ),
	.delay_reg_1_3(\delay_line_inst|delay_reg[3][1]~q ),
	.delay_reg_2_3(\delay_line_inst|delay_reg[3][2]~q ),
	.delay_reg_3_3(\delay_line_inst|delay_reg[3][3]~q ),
	.delay_reg_4_3(\delay_line_inst|delay_reg[3][4]~q ),
	.delay_reg_5_3(\delay_line_inst|delay_reg[3][5]~q ),
	.delay_reg_6_3(\delay_line_inst|delay_reg[3][6]~q ),
	.delay_reg_7_3(\delay_line_inst|delay_reg[3][7]~q ),
	.delay_reg_8_3(\delay_line_inst|delay_reg[3][8]~q ),
	.delay_reg_9_3(\delay_line_inst|delay_reg[3][9]~q ),
	.delay_reg_10_3(\delay_line_inst|delay_reg[3][10]~q ),
	.delay_reg_11_3(\delay_line_inst|delay_reg[3][11]~q ),
	.delay_reg_12_3(\delay_line_inst|delay_reg[3][12]~q ),
	.delay_reg_13_3(\delay_line_inst|delay_reg[3][13]~q ),
	.delay_reg_14_3(\delay_line_inst|delay_reg[3][14]~q ),
	.delay_reg_15_3(\delay_line_inst|delay_reg[3][15]~q ),
	.delay_reg_16_3(\delay_line_inst|delay_reg[3][16]~q ),
	.delay_reg_17_3(\delay_line_inst|delay_reg[3][17]~q ),
	.delay_reg_18_3(\delay_line_inst|delay_reg[3][18]~q ),
	.delay_reg_19_3(\delay_line_inst|delay_reg[3][19]~q ),
	.delay_reg_20_3(\delay_line_inst|delay_reg[3][20]~q ),
	.delay_reg_21_3(\delay_line_inst|delay_reg[3][21]~q ),
	.delay_reg_22_3(\delay_line_inst|delay_reg[3][22]~q ),
	.delay_reg_23_3(\delay_line_inst|delay_reg[3][23]~q ),
	.delay_reg_24_3(delay_reg_24_3),
	.clock(clk_clk),
	.ppd_cfg_enable(ppd_cfg_enable));

fiftyfivenm_lcell_comb \avalon_streaming_source_data[0]~1 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_0),
	.cout());
defparam \avalon_streaming_source_data[0]~1 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[1]~2 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_1),
	.cout());
defparam \avalon_streaming_source_data[1]~2 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[1]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[2]~3 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_2),
	.cout());
defparam \avalon_streaming_source_data[2]~3 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[2]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[3]~4 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_3),
	.cout());
defparam \avalon_streaming_source_data[3]~4 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[3]~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[4]~5 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_4),
	.cout());
defparam \avalon_streaming_source_data[4]~5 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[4]~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[5]~6 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_5),
	.cout());
defparam \avalon_streaming_source_data[5]~6 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[5]~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[6]~7 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_6),
	.cout());
defparam \avalon_streaming_source_data[6]~7 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[6]~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[7]~8 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_7),
	.cout());
defparam \avalon_streaming_source_data[7]~8 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[7]~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[8]~9 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_8),
	.cout());
defparam \avalon_streaming_source_data[8]~9 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[8]~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[9]~10 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_9),
	.cout());
defparam \avalon_streaming_source_data[9]~10 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[9]~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[10]~11 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_10),
	.cout());
defparam \avalon_streaming_source_data[10]~11 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[10]~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[11]~12 (
	.dataa(\delay_line_inst|delay_reg[3][11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avalon_streaming_source_data~0_combout ),
	.cin(gnd),
	.combout(avalon_streaming_source_data_11),
	.cout());
defparam \avalon_streaming_source_data[11]~12 .lut_mask = 16'h00AA;
defparam \avalon_streaming_source_data[11]~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[12]~13 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_12),
	.cout());
defparam \avalon_streaming_source_data[12]~13 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[12]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[13]~14 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_13),
	.cout());
defparam \avalon_streaming_source_data[13]~14 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[13]~14 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[14]~15 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_14),
	.cout());
defparam \avalon_streaming_source_data[14]~15 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[14]~15 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[15]~16 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_15),
	.cout());
defparam \avalon_streaming_source_data[15]~16 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[15]~16 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[16]~17 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_16),
	.cout());
defparam \avalon_streaming_source_data[16]~17 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[16]~17 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[17]~18 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][17]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_17),
	.cout());
defparam \avalon_streaming_source_data[17]~18 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[17]~18 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[18]~19 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][18]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_18),
	.cout());
defparam \avalon_streaming_source_data[18]~19 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[18]~19 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[19]~20 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][19]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_19),
	.cout());
defparam \avalon_streaming_source_data[19]~20 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[19]~20 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[20]~21 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_20),
	.cout());
defparam \avalon_streaming_source_data[20]~21 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[20]~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[21]~22 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][21]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_21),
	.cout());
defparam \avalon_streaming_source_data[21]~22 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[21]~22 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[22]~23 (
	.dataa(\avalon_streaming_source_data~0_combout ),
	.datab(\delay_line_inst|delay_reg[3][22]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(avalon_streaming_source_data_22),
	.cout());
defparam \avalon_streaming_source_data[22]~23 .lut_mask = 16'hEEEE;
defparam \avalon_streaming_source_data[22]~23 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data[23]~24 (
	.dataa(\delay_line_inst|delay_reg[3][23]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avalon_streaming_source_data~0_combout ),
	.cin(gnd),
	.combout(avalon_streaming_source_data_23),
	.cout());
defparam \avalon_streaming_source_data[23]~24 .lut_mask = 16'h00AA;
defparam \avalon_streaming_source_data[23]~24 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \avalon_streaming_source_data~0 (
	.dataa(\running_sum_inst|LessThan0~34_combout ),
	.datab(\running_sum_inst|launch~2_combout ),
	.datac(\delay_line_inst|delay_reg[2][25]~q ),
	.datad(\running_sum_inst|long_shift_rescale[25]~q ),
	.cin(gnd),
	.combout(\avalon_streaming_source_data~0_combout ),
	.cout());
defparam \avalon_streaming_source_data~0 .lut_mask = 16'h0080;
defparam \avalon_streaming_source_data~0 .sum_lutc_input = "datac";

endmodule

module lms_dsp_cmplx2mag (
	mag_reg_0,
	mag_reg_1,
	mag_reg_2,
	mag_reg_3,
	mag_reg_4,
	mag_reg_5,
	mag_reg_6,
	mag_reg_7,
	mag_reg_8,
	mag_reg_9,
	mag_reg_10,
	mag_reg_11,
	mag_reg_12,
	altera_reset_synchronizer_int_chain_out,
	data_out_12,
	data_out_0,
	data_out_11,
	data_out_10,
	data_out_9,
	data_out_8,
	data_out_7,
	data_out_6,
	data_out_5,
	data_out_4,
	data_out_3,
	data_out_2,
	data_out_1,
	data_out_23,
	data_out_22,
	data_out_21,
	data_out_20,
	data_out_19,
	data_out_18,
	data_out_17,
	data_out_16,
	data_out_15,
	data_out_14,
	data_out_13,
	clock)/* synthesis synthesis_greybox=0 */;
output 	mag_reg_0;
output 	mag_reg_1;
output 	mag_reg_2;
output 	mag_reg_3;
output 	mag_reg_4;
output 	mag_reg_5;
output 	mag_reg_6;
output 	mag_reg_7;
output 	mag_reg_8;
output 	mag_reg_9;
output 	mag_reg_10;
output 	mag_reg_11;
output 	mag_reg_12;
input 	altera_reset_synchronizer_int_chain_out;
input 	data_out_12;
input 	data_out_0;
input 	data_out_11;
input 	data_out_10;
input 	data_out_9;
input 	data_out_8;
input 	data_out_7;
input 	data_out_6;
input 	data_out_5;
input 	data_out_4;
input 	data_out_3;
input 	data_out_2;
input 	data_out_1;
input 	data_out_23;
input 	data_out_22;
input 	data_out_21;
input 	data_out_20;
input 	data_out_19;
input 	data_out_18;
input 	data_out_17;
input 	data_out_16;
input 	data_out_15;
input 	data_out_14;
input 	data_out_13;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add1~1_cout ;
wire \Add1~3 ;
wire \Add1~5 ;
wire \Add1~7 ;
wire \Add1~9 ;
wire \Add1~11 ;
wire \Add1~13 ;
wire \Add1~15 ;
wire \Add1~17 ;
wire \Add1~19 ;
wire \Add1~21 ;
wire \Add1~22_combout ;
wire \abs_q[11]~0_combout ;
wire \Add0~1_cout ;
wire \Add0~3 ;
wire \Add0~5 ;
wire \Add0~7 ;
wire \Add0~9 ;
wire \Add0~11 ;
wire \Add0~13 ;
wire \Add0~15 ;
wire \Add0~17 ;
wire \Add0~19 ;
wire \Add0~21 ;
wire \Add0~22_combout ;
wire \abs_i[11]~0_combout ;
wire \Add1~20_combout ;
wire \abs_q[10]~1_combout ;
wire \Add0~20_combout ;
wire \abs_i[10]~1_combout ;
wire \Add1~18_combout ;
wire \abs_q[9]~2_combout ;
wire \Add0~18_combout ;
wire \abs_i[9]~2_combout ;
wire \Add1~16_combout ;
wire \abs_q[8]~3_combout ;
wire \Add0~16_combout ;
wire \abs_i[8]~3_combout ;
wire \Add1~14_combout ;
wire \abs_q[7]~4_combout ;
wire \Add0~14_combout ;
wire \abs_i[7]~4_combout ;
wire \Add1~12_combout ;
wire \abs_q[6]~5_combout ;
wire \Add0~12_combout ;
wire \abs_i[6]~5_combout ;
wire \Add1~10_combout ;
wire \abs_q[5]~6_combout ;
wire \Add0~10_combout ;
wire \abs_i[5]~6_combout ;
wire \Add1~8_combout ;
wire \abs_q[4]~7_combout ;
wire \Add0~8_combout ;
wire \abs_i[4]~7_combout ;
wire \Add1~6_combout ;
wire \abs_q[3]~8_combout ;
wire \Add0~6_combout ;
wire \abs_i[3]~8_combout ;
wire \Add1~4_combout ;
wire \abs_q[2]~9_combout ;
wire \Add0~4_combout ;
wire \abs_i[2]~9_combout ;
wire \Add1~2_combout ;
wire \abs_q[1]~10_combout ;
wire \Add0~2_combout ;
wire \abs_i[1]~10_combout ;
wire \LessThan0~1_cout ;
wire \LessThan0~3_cout ;
wire \LessThan0~5_cout ;
wire \LessThan0~7_cout ;
wire \LessThan0~9_cout ;
wire \LessThan0~11_cout ;
wire \LessThan0~13_cout ;
wire \LessThan0~15_cout ;
wire \LessThan0~17_cout ;
wire \LessThan0~19_cout ;
wire \LessThan0~21_cout ;
wire \LessThan0~22_combout ;
wire \max[0]~0_combout ;
wire \min[2]~4_combout ;
wire \mag_reg[0]~13_combout ;
wire \max[1]~1_combout ;
wire \min[3]~5_combout ;
wire \mag_reg[0]~14 ;
wire \mag_reg[1]~15_combout ;
wire \max[2]~2_combout ;
wire \min[4]~6_combout ;
wire \mag_reg[1]~16 ;
wire \mag_reg[2]~17_combout ;
wire \max[3]~3_combout ;
wire \min[5]~7_combout ;
wire \mag_reg[2]~18 ;
wire \mag_reg[3]~19_combout ;
wire \max[4]~4_combout ;
wire \min[6]~8_combout ;
wire \mag_reg[3]~20 ;
wire \mag_reg[4]~21_combout ;
wire \max[5]~5_combout ;
wire \min[7]~9_combout ;
wire \mag_reg[4]~22 ;
wire \mag_reg[5]~23_combout ;
wire \max[6]~6_combout ;
wire \min[8]~10_combout ;
wire \mag_reg[5]~24 ;
wire \mag_reg[6]~25_combout ;
wire \max[7]~7_combout ;
wire \min[9]~11_combout ;
wire \mag_reg[6]~26 ;
wire \mag_reg[7]~27_combout ;
wire \max[8]~8_combout ;
wire \min[10]~12_combout ;
wire \mag_reg[7]~28 ;
wire \mag_reg[8]~29_combout ;
wire \min[11]~13_combout ;
wire \max[9]~9_combout ;
wire \mag_reg[8]~30 ;
wire \mag_reg[9]~31_combout ;
wire \max[10]~10_combout ;
wire \mag_reg[9]~32 ;
wire \mag_reg[10]~33_combout ;
wire \max[11]~11_combout ;
wire \max[11]~12_combout ;
wire \mag_reg[10]~34 ;
wire \mag_reg[11]~35_combout ;
wire \mag_reg[11]~36 ;
wire \mag_reg[12]~37_combout ;


dffeas \mag_reg[0] (
	.clk(clock),
	.d(\mag_reg[0]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(mag_reg_0),
	.prn(vcc));
defparam \mag_reg[0] .is_wysiwyg = "true";
defparam \mag_reg[0] .power_up = "low";

dffeas \mag_reg[1] (
	.clk(clock),
	.d(\mag_reg[1]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(mag_reg_1),
	.prn(vcc));
defparam \mag_reg[1] .is_wysiwyg = "true";
defparam \mag_reg[1] .power_up = "low";

dffeas \mag_reg[2] (
	.clk(clock),
	.d(\mag_reg[2]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(mag_reg_2),
	.prn(vcc));
defparam \mag_reg[2] .is_wysiwyg = "true";
defparam \mag_reg[2] .power_up = "low";

dffeas \mag_reg[3] (
	.clk(clock),
	.d(\mag_reg[3]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(mag_reg_3),
	.prn(vcc));
defparam \mag_reg[3] .is_wysiwyg = "true";
defparam \mag_reg[3] .power_up = "low";

dffeas \mag_reg[4] (
	.clk(clock),
	.d(\mag_reg[4]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(mag_reg_4),
	.prn(vcc));
defparam \mag_reg[4] .is_wysiwyg = "true";
defparam \mag_reg[4] .power_up = "low";

dffeas \mag_reg[5] (
	.clk(clock),
	.d(\mag_reg[5]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(mag_reg_5),
	.prn(vcc));
defparam \mag_reg[5] .is_wysiwyg = "true";
defparam \mag_reg[5] .power_up = "low";

dffeas \mag_reg[6] (
	.clk(clock),
	.d(\mag_reg[6]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(mag_reg_6),
	.prn(vcc));
defparam \mag_reg[6] .is_wysiwyg = "true";
defparam \mag_reg[6] .power_up = "low";

dffeas \mag_reg[7] (
	.clk(clock),
	.d(\mag_reg[7]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(mag_reg_7),
	.prn(vcc));
defparam \mag_reg[7] .is_wysiwyg = "true";
defparam \mag_reg[7] .power_up = "low";

dffeas \mag_reg[8] (
	.clk(clock),
	.d(\mag_reg[8]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(mag_reg_8),
	.prn(vcc));
defparam \mag_reg[8] .is_wysiwyg = "true";
defparam \mag_reg[8] .power_up = "low";

dffeas \mag_reg[9] (
	.clk(clock),
	.d(\mag_reg[9]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(mag_reg_9),
	.prn(vcc));
defparam \mag_reg[9] .is_wysiwyg = "true";
defparam \mag_reg[9] .power_up = "low";

dffeas \mag_reg[10] (
	.clk(clock),
	.d(\mag_reg[10]~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(mag_reg_10),
	.prn(vcc));
defparam \mag_reg[10] .is_wysiwyg = "true";
defparam \mag_reg[10] .power_up = "low";

dffeas \mag_reg[11] (
	.clk(clock),
	.d(\mag_reg[11]~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(mag_reg_11),
	.prn(vcc));
defparam \mag_reg[11] .is_wysiwyg = "true";
defparam \mag_reg[11] .power_up = "low";

dffeas \mag_reg[12] (
	.clk(clock),
	.d(\mag_reg[12]~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(mag_reg_12),
	.prn(vcc));
defparam \mag_reg[12] .is_wysiwyg = "true";
defparam \mag_reg[12] .power_up = "low";

fiftyfivenm_lcell_comb \Add1~1 (
	.dataa(data_out_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\Add1~1_cout ));
defparam \Add1~1 .lut_mask = 16'h0055;
defparam \Add1~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add1~2 (
	.dataa(data_out_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1_cout ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
defparam \Add1~2 .lut_mask = 16'hA5AF;
defparam \Add1~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add1~4 (
	.dataa(data_out_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
defparam \Add1~4 .lut_mask = 16'h5A05;
defparam \Add1~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add1~6 (
	.dataa(data_out_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
defparam \Add1~6 .lut_mask = 16'hA5AF;
defparam \Add1~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add1~8 (
	.dataa(data_out_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
defparam \Add1~8 .lut_mask = 16'h5A05;
defparam \Add1~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add1~10 (
	.dataa(data_out_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout(\Add1~11 ));
defparam \Add1~10 .lut_mask = 16'hA5AF;
defparam \Add1~10 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add1~12 (
	.dataa(data_out_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~11 ),
	.combout(\Add1~12_combout ),
	.cout(\Add1~13 ));
defparam \Add1~12 .lut_mask = 16'h5A05;
defparam \Add1~12 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add1~14 (
	.dataa(data_out_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~13 ),
	.combout(\Add1~14_combout ),
	.cout(\Add1~15 ));
defparam \Add1~14 .lut_mask = 16'hA5AF;
defparam \Add1~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add1~16 (
	.dataa(data_out_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~15 ),
	.combout(\Add1~16_combout ),
	.cout(\Add1~17 ));
defparam \Add1~16 .lut_mask = 16'h5A05;
defparam \Add1~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add1~18 (
	.dataa(data_out_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~17 ),
	.combout(\Add1~18_combout ),
	.cout(\Add1~19 ));
defparam \Add1~18 .lut_mask = 16'hA5AF;
defparam \Add1~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add1~20 (
	.dataa(data_out_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~19 ),
	.combout(\Add1~20_combout ),
	.cout(\Add1~21 ));
defparam \Add1~20 .lut_mask = 16'h5A05;
defparam \Add1~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add1~22 (
	.dataa(data_out_11),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add1~21 ),
	.combout(\Add1~22_combout ),
	.cout());
defparam \Add1~22 .lut_mask = 16'hA5A5;
defparam \Add1~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \abs_q[11]~0 (
	.dataa(data_out_11),
	.datab(\Add1~22_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\abs_q[11]~0_combout ),
	.cout());
defparam \abs_q[11]~0 .lut_mask = 16'h8888;
defparam \abs_q[11]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~1 (
	.dataa(data_out_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\Add0~1_cout ));
defparam \Add0~1 .lut_mask = 16'h0055;
defparam \Add0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~2 (
	.dataa(data_out_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1_cout ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'hA5AF;
defparam \Add0~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~4 (
	.dataa(data_out_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'h5A05;
defparam \Add0~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~6 (
	.dataa(data_out_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'hA5AF;
defparam \Add0~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~8 (
	.dataa(data_out_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
defparam \Add0~8 .lut_mask = 16'h5A05;
defparam \Add0~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~10 (
	.dataa(data_out_17),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
defparam \Add0~10 .lut_mask = 16'hA5AF;
defparam \Add0~10 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~12 (
	.dataa(data_out_18),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
defparam \Add0~12 .lut_mask = 16'h5A05;
defparam \Add0~12 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~14 (
	.dataa(data_out_19),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
defparam \Add0~14 .lut_mask = 16'hA5AF;
defparam \Add0~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~16 (
	.dataa(data_out_20),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout(\Add0~17 ));
defparam \Add0~16 .lut_mask = 16'h5A05;
defparam \Add0~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~18 (
	.dataa(data_out_21),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~17 ),
	.combout(\Add0~18_combout ),
	.cout(\Add0~19 ));
defparam \Add0~18 .lut_mask = 16'hA5AF;
defparam \Add0~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~20 (
	.dataa(data_out_22),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~19 ),
	.combout(\Add0~20_combout ),
	.cout(\Add0~21 ));
defparam \Add0~20 .lut_mask = 16'h5A05;
defparam \Add0~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~22 (
	.dataa(data_out_23),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~21 ),
	.combout(\Add0~22_combout ),
	.cout());
defparam \Add0~22 .lut_mask = 16'hA5A5;
defparam \Add0~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \abs_i[11]~0 (
	.dataa(data_out_23),
	.datab(\Add0~22_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\abs_i[11]~0_combout ),
	.cout());
defparam \abs_i[11]~0 .lut_mask = 16'h8888;
defparam \abs_i[11]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_q[10]~1 (
	.dataa(\Add1~20_combout ),
	.datab(data_out_10),
	.datac(gnd),
	.datad(data_out_11),
	.cin(gnd),
	.combout(\abs_q[10]~1_combout ),
	.cout());
defparam \abs_q[10]~1 .lut_mask = 16'hAACC;
defparam \abs_q[10]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_i[10]~1 (
	.dataa(\Add0~20_combout ),
	.datab(data_out_22),
	.datac(gnd),
	.datad(data_out_23),
	.cin(gnd),
	.combout(\abs_i[10]~1_combout ),
	.cout());
defparam \abs_i[10]~1 .lut_mask = 16'hAACC;
defparam \abs_i[10]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_q[9]~2 (
	.dataa(\Add1~18_combout ),
	.datab(data_out_9),
	.datac(gnd),
	.datad(data_out_11),
	.cin(gnd),
	.combout(\abs_q[9]~2_combout ),
	.cout());
defparam \abs_q[9]~2 .lut_mask = 16'hAACC;
defparam \abs_q[9]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_i[9]~2 (
	.dataa(\Add0~18_combout ),
	.datab(data_out_21),
	.datac(gnd),
	.datad(data_out_23),
	.cin(gnd),
	.combout(\abs_i[9]~2_combout ),
	.cout());
defparam \abs_i[9]~2 .lut_mask = 16'hAACC;
defparam \abs_i[9]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_q[8]~3 (
	.dataa(\Add1~16_combout ),
	.datab(data_out_8),
	.datac(gnd),
	.datad(data_out_11),
	.cin(gnd),
	.combout(\abs_q[8]~3_combout ),
	.cout());
defparam \abs_q[8]~3 .lut_mask = 16'hAACC;
defparam \abs_q[8]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_i[8]~3 (
	.dataa(\Add0~16_combout ),
	.datab(data_out_20),
	.datac(gnd),
	.datad(data_out_23),
	.cin(gnd),
	.combout(\abs_i[8]~3_combout ),
	.cout());
defparam \abs_i[8]~3 .lut_mask = 16'hAACC;
defparam \abs_i[8]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_q[7]~4 (
	.dataa(\Add1~14_combout ),
	.datab(data_out_7),
	.datac(gnd),
	.datad(data_out_11),
	.cin(gnd),
	.combout(\abs_q[7]~4_combout ),
	.cout());
defparam \abs_q[7]~4 .lut_mask = 16'hAACC;
defparam \abs_q[7]~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_i[7]~4 (
	.dataa(\Add0~14_combout ),
	.datab(data_out_19),
	.datac(gnd),
	.datad(data_out_23),
	.cin(gnd),
	.combout(\abs_i[7]~4_combout ),
	.cout());
defparam \abs_i[7]~4 .lut_mask = 16'hAACC;
defparam \abs_i[7]~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_q[6]~5 (
	.dataa(\Add1~12_combout ),
	.datab(data_out_6),
	.datac(gnd),
	.datad(data_out_11),
	.cin(gnd),
	.combout(\abs_q[6]~5_combout ),
	.cout());
defparam \abs_q[6]~5 .lut_mask = 16'hAACC;
defparam \abs_q[6]~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_i[6]~5 (
	.dataa(\Add0~12_combout ),
	.datab(data_out_18),
	.datac(gnd),
	.datad(data_out_23),
	.cin(gnd),
	.combout(\abs_i[6]~5_combout ),
	.cout());
defparam \abs_i[6]~5 .lut_mask = 16'hAACC;
defparam \abs_i[6]~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_q[5]~6 (
	.dataa(\Add1~10_combout ),
	.datab(data_out_5),
	.datac(gnd),
	.datad(data_out_11),
	.cin(gnd),
	.combout(\abs_q[5]~6_combout ),
	.cout());
defparam \abs_q[5]~6 .lut_mask = 16'hAACC;
defparam \abs_q[5]~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_i[5]~6 (
	.dataa(\Add0~10_combout ),
	.datab(data_out_17),
	.datac(gnd),
	.datad(data_out_23),
	.cin(gnd),
	.combout(\abs_i[5]~6_combout ),
	.cout());
defparam \abs_i[5]~6 .lut_mask = 16'hAACC;
defparam \abs_i[5]~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_q[4]~7 (
	.dataa(\Add1~8_combout ),
	.datab(data_out_4),
	.datac(gnd),
	.datad(data_out_11),
	.cin(gnd),
	.combout(\abs_q[4]~7_combout ),
	.cout());
defparam \abs_q[4]~7 .lut_mask = 16'hAACC;
defparam \abs_q[4]~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_i[4]~7 (
	.dataa(\Add0~8_combout ),
	.datab(data_out_16),
	.datac(gnd),
	.datad(data_out_23),
	.cin(gnd),
	.combout(\abs_i[4]~7_combout ),
	.cout());
defparam \abs_i[4]~7 .lut_mask = 16'hAACC;
defparam \abs_i[4]~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_q[3]~8 (
	.dataa(\Add1~6_combout ),
	.datab(data_out_3),
	.datac(gnd),
	.datad(data_out_11),
	.cin(gnd),
	.combout(\abs_q[3]~8_combout ),
	.cout());
defparam \abs_q[3]~8 .lut_mask = 16'hAACC;
defparam \abs_q[3]~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_i[3]~8 (
	.dataa(\Add0~6_combout ),
	.datab(data_out_15),
	.datac(gnd),
	.datad(data_out_23),
	.cin(gnd),
	.combout(\abs_i[3]~8_combout ),
	.cout());
defparam \abs_i[3]~8 .lut_mask = 16'hAACC;
defparam \abs_i[3]~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_q[2]~9 (
	.dataa(\Add1~4_combout ),
	.datab(data_out_2),
	.datac(gnd),
	.datad(data_out_11),
	.cin(gnd),
	.combout(\abs_q[2]~9_combout ),
	.cout());
defparam \abs_q[2]~9 .lut_mask = 16'hAACC;
defparam \abs_q[2]~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_i[2]~9 (
	.dataa(\Add0~4_combout ),
	.datab(data_out_14),
	.datac(gnd),
	.datad(data_out_23),
	.cin(gnd),
	.combout(\abs_i[2]~9_combout ),
	.cout());
defparam \abs_i[2]~9 .lut_mask = 16'hAACC;
defparam \abs_i[2]~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_q[1]~10 (
	.dataa(\Add1~2_combout ),
	.datab(data_out_1),
	.datac(gnd),
	.datad(data_out_11),
	.cin(gnd),
	.combout(\abs_q[1]~10_combout ),
	.cout());
defparam \abs_q[1]~10 .lut_mask = 16'hAACC;
defparam \abs_q[1]~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \abs_i[1]~10 (
	.dataa(\Add0~2_combout ),
	.datab(data_out_13),
	.datac(gnd),
	.datad(data_out_23),
	.cin(gnd),
	.combout(\abs_i[1]~10_combout ),
	.cout());
defparam \abs_i[1]~10 .lut_mask = 16'hAACC;
defparam \abs_i[1]~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \LessThan0~1 (
	.dataa(data_out_0),
	.datab(data_out_12),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan0~1_cout ));
defparam \LessThan0~1 .lut_mask = 16'h0044;
defparam \LessThan0~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~3 (
	.dataa(\abs_q[1]~10_combout ),
	.datab(\abs_i[1]~10_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~1_cout ),
	.combout(),
	.cout(\LessThan0~3_cout ));
defparam \LessThan0~3 .lut_mask = 16'h002B;
defparam \LessThan0~3 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~5 (
	.dataa(\abs_q[2]~9_combout ),
	.datab(\abs_i[2]~9_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~3_cout ),
	.combout(),
	.cout(\LessThan0~5_cout ));
defparam \LessThan0~5 .lut_mask = 16'h004D;
defparam \LessThan0~5 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~7 (
	.dataa(\abs_q[3]~8_combout ),
	.datab(\abs_i[3]~8_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~5_cout ),
	.combout(),
	.cout(\LessThan0~7_cout ));
defparam \LessThan0~7 .lut_mask = 16'h002B;
defparam \LessThan0~7 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~9 (
	.dataa(\abs_q[4]~7_combout ),
	.datab(\abs_i[4]~7_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~7_cout ),
	.combout(),
	.cout(\LessThan0~9_cout ));
defparam \LessThan0~9 .lut_mask = 16'h004D;
defparam \LessThan0~9 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~11 (
	.dataa(\abs_q[5]~6_combout ),
	.datab(\abs_i[5]~6_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~9_cout ),
	.combout(),
	.cout(\LessThan0~11_cout ));
defparam \LessThan0~11 .lut_mask = 16'h002B;
defparam \LessThan0~11 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~13 (
	.dataa(\abs_q[6]~5_combout ),
	.datab(\abs_i[6]~5_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~11_cout ),
	.combout(),
	.cout(\LessThan0~13_cout ));
defparam \LessThan0~13 .lut_mask = 16'h004D;
defparam \LessThan0~13 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~15 (
	.dataa(\abs_q[7]~4_combout ),
	.datab(\abs_i[7]~4_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~13_cout ),
	.combout(),
	.cout(\LessThan0~15_cout ));
defparam \LessThan0~15 .lut_mask = 16'h002B;
defparam \LessThan0~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~17 (
	.dataa(\abs_q[8]~3_combout ),
	.datab(\abs_i[8]~3_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~15_cout ),
	.combout(),
	.cout(\LessThan0~17_cout ));
defparam \LessThan0~17 .lut_mask = 16'h004D;
defparam \LessThan0~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~19 (
	.dataa(\abs_q[9]~2_combout ),
	.datab(\abs_i[9]~2_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~17_cout ),
	.combout(),
	.cout(\LessThan0~19_cout ));
defparam \LessThan0~19 .lut_mask = 16'h002B;
defparam \LessThan0~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~21 (
	.dataa(\abs_q[10]~1_combout ),
	.datab(\abs_i[10]~1_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~19_cout ),
	.combout(),
	.cout(\LessThan0~21_cout ));
defparam \LessThan0~21 .lut_mask = 16'h004D;
defparam \LessThan0~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~22 (
	.dataa(\abs_q[11]~0_combout ),
	.datab(\abs_i[11]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(\LessThan0~21_cout ),
	.combout(\LessThan0~22_combout ),
	.cout());
defparam \LessThan0~22 .lut_mask = 16'hD4D4;
defparam \LessThan0~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \max[0]~0 (
	.dataa(data_out_12),
	.datab(data_out_0),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\max[0]~0_combout ),
	.cout());
defparam \max[0]~0 .lut_mask = 16'hAACC;
defparam \max[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \min[2]~4 (
	.dataa(\abs_q[2]~9_combout ),
	.datab(\abs_i[2]~9_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\min[2]~4_combout ),
	.cout());
defparam \min[2]~4 .lut_mask = 16'hAACC;
defparam \min[2]~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mag_reg[0]~13 (
	.dataa(\max[0]~0_combout ),
	.datab(\min[2]~4_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\mag_reg[0]~13_combout ),
	.cout(\mag_reg[0]~14 ));
defparam \mag_reg[0]~13 .lut_mask = 16'h6688;
defparam \mag_reg[0]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \max[1]~1 (
	.dataa(\abs_i[1]~10_combout ),
	.datab(\abs_q[1]~10_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\max[1]~1_combout ),
	.cout());
defparam \max[1]~1 .lut_mask = 16'hAACC;
defparam \max[1]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \min[3]~5 (
	.dataa(\abs_q[3]~8_combout ),
	.datab(\abs_i[3]~8_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\min[3]~5_combout ),
	.cout());
defparam \min[3]~5 .lut_mask = 16'hAACC;
defparam \min[3]~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mag_reg[1]~15 (
	.dataa(\max[1]~1_combout ),
	.datab(\min[3]~5_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\mag_reg[0]~14 ),
	.combout(\mag_reg[1]~15_combout ),
	.cout(\mag_reg[1]~16 ));
defparam \mag_reg[1]~15 .lut_mask = 16'h9617;
defparam \mag_reg[1]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \max[2]~2 (
	.dataa(\abs_i[2]~9_combout ),
	.datab(\abs_q[2]~9_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\max[2]~2_combout ),
	.cout());
defparam \max[2]~2 .lut_mask = 16'hAACC;
defparam \max[2]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \min[4]~6 (
	.dataa(\abs_q[4]~7_combout ),
	.datab(\abs_i[4]~7_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\min[4]~6_combout ),
	.cout());
defparam \min[4]~6 .lut_mask = 16'hAACC;
defparam \min[4]~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mag_reg[2]~17 (
	.dataa(\max[2]~2_combout ),
	.datab(\min[4]~6_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\mag_reg[1]~16 ),
	.combout(\mag_reg[2]~17_combout ),
	.cout(\mag_reg[2]~18 ));
defparam \mag_reg[2]~17 .lut_mask = 16'h698E;
defparam \mag_reg[2]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \max[3]~3 (
	.dataa(\abs_i[3]~8_combout ),
	.datab(\abs_q[3]~8_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\max[3]~3_combout ),
	.cout());
defparam \max[3]~3 .lut_mask = 16'hAACC;
defparam \max[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \min[5]~7 (
	.dataa(\abs_q[5]~6_combout ),
	.datab(\abs_i[5]~6_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\min[5]~7_combout ),
	.cout());
defparam \min[5]~7 .lut_mask = 16'hAACC;
defparam \min[5]~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mag_reg[3]~19 (
	.dataa(\max[3]~3_combout ),
	.datab(\min[5]~7_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\mag_reg[2]~18 ),
	.combout(\mag_reg[3]~19_combout ),
	.cout(\mag_reg[3]~20 ));
defparam \mag_reg[3]~19 .lut_mask = 16'h9617;
defparam \mag_reg[3]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \max[4]~4 (
	.dataa(\abs_i[4]~7_combout ),
	.datab(\abs_q[4]~7_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\max[4]~4_combout ),
	.cout());
defparam \max[4]~4 .lut_mask = 16'hAACC;
defparam \max[4]~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \min[6]~8 (
	.dataa(\abs_q[6]~5_combout ),
	.datab(\abs_i[6]~5_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\min[6]~8_combout ),
	.cout());
defparam \min[6]~8 .lut_mask = 16'hAACC;
defparam \min[6]~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mag_reg[4]~21 (
	.dataa(\max[4]~4_combout ),
	.datab(\min[6]~8_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\mag_reg[3]~20 ),
	.combout(\mag_reg[4]~21_combout ),
	.cout(\mag_reg[4]~22 ));
defparam \mag_reg[4]~21 .lut_mask = 16'h698E;
defparam \mag_reg[4]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \max[5]~5 (
	.dataa(\abs_i[5]~6_combout ),
	.datab(\abs_q[5]~6_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\max[5]~5_combout ),
	.cout());
defparam \max[5]~5 .lut_mask = 16'hAACC;
defparam \max[5]~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \min[7]~9 (
	.dataa(\abs_q[7]~4_combout ),
	.datab(\abs_i[7]~4_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\min[7]~9_combout ),
	.cout());
defparam \min[7]~9 .lut_mask = 16'hAACC;
defparam \min[7]~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mag_reg[5]~23 (
	.dataa(\max[5]~5_combout ),
	.datab(\min[7]~9_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\mag_reg[4]~22 ),
	.combout(\mag_reg[5]~23_combout ),
	.cout(\mag_reg[5]~24 ));
defparam \mag_reg[5]~23 .lut_mask = 16'h9617;
defparam \mag_reg[5]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \max[6]~6 (
	.dataa(\abs_i[6]~5_combout ),
	.datab(\abs_q[6]~5_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\max[6]~6_combout ),
	.cout());
defparam \max[6]~6 .lut_mask = 16'hAACC;
defparam \max[6]~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \min[8]~10 (
	.dataa(\abs_q[8]~3_combout ),
	.datab(\abs_i[8]~3_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\min[8]~10_combout ),
	.cout());
defparam \min[8]~10 .lut_mask = 16'hAACC;
defparam \min[8]~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mag_reg[6]~25 (
	.dataa(\max[6]~6_combout ),
	.datab(\min[8]~10_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\mag_reg[5]~24 ),
	.combout(\mag_reg[6]~25_combout ),
	.cout(\mag_reg[6]~26 ));
defparam \mag_reg[6]~25 .lut_mask = 16'h698E;
defparam \mag_reg[6]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \max[7]~7 (
	.dataa(\abs_i[7]~4_combout ),
	.datab(\abs_q[7]~4_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\max[7]~7_combout ),
	.cout());
defparam \max[7]~7 .lut_mask = 16'hAACC;
defparam \max[7]~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \min[9]~11 (
	.dataa(\abs_q[9]~2_combout ),
	.datab(\abs_i[9]~2_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\min[9]~11_combout ),
	.cout());
defparam \min[9]~11 .lut_mask = 16'hAACC;
defparam \min[9]~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mag_reg[7]~27 (
	.dataa(\max[7]~7_combout ),
	.datab(\min[9]~11_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\mag_reg[6]~26 ),
	.combout(\mag_reg[7]~27_combout ),
	.cout(\mag_reg[7]~28 ));
defparam \mag_reg[7]~27 .lut_mask = 16'h9617;
defparam \mag_reg[7]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \max[8]~8 (
	.dataa(\abs_i[8]~3_combout ),
	.datab(\abs_q[8]~3_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\max[8]~8_combout ),
	.cout());
defparam \max[8]~8 .lut_mask = 16'hAACC;
defparam \max[8]~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \min[10]~12 (
	.dataa(\abs_q[10]~1_combout ),
	.datab(\abs_i[10]~1_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\min[10]~12_combout ),
	.cout());
defparam \min[10]~12 .lut_mask = 16'hAACC;
defparam \min[10]~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mag_reg[8]~29 (
	.dataa(\max[8]~8_combout ),
	.datab(\min[10]~12_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\mag_reg[7]~28 ),
	.combout(\mag_reg[8]~29_combout ),
	.cout(\mag_reg[8]~30 ));
defparam \mag_reg[8]~29 .lut_mask = 16'h698E;
defparam \mag_reg[8]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \min[11]~13 (
	.dataa(data_out_11),
	.datab(\Add1~22_combout ),
	.datac(\abs_i[11]~0_combout ),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\min[11]~13_combout ),
	.cout());
defparam \min[11]~13 .lut_mask = 16'h88F0;
defparam \min[11]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \max[9]~9 (
	.dataa(\abs_i[9]~2_combout ),
	.datab(\abs_q[9]~2_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\max[9]~9_combout ),
	.cout());
defparam \max[9]~9 .lut_mask = 16'hAACC;
defparam \max[9]~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mag_reg[9]~31 (
	.dataa(\min[11]~13_combout ),
	.datab(\max[9]~9_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\mag_reg[8]~30 ),
	.combout(\mag_reg[9]~31_combout ),
	.cout(\mag_reg[9]~32 ));
defparam \mag_reg[9]~31 .lut_mask = 16'h9617;
defparam \mag_reg[9]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \max[10]~10 (
	.dataa(\abs_i[10]~1_combout ),
	.datab(\abs_q[10]~1_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\max[10]~10_combout ),
	.cout());
defparam \max[10]~10 .lut_mask = 16'hAACC;
defparam \max[10]~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mag_reg[10]~33 (
	.dataa(\max[10]~10_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\mag_reg[9]~32 ),
	.combout(\mag_reg[10]~33_combout ),
	.cout(\mag_reg[10]~34 ));
defparam \mag_reg[10]~33 .lut_mask = 16'hA50A;
defparam \mag_reg[10]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \max[11]~11 (
	.dataa(data_out_23),
	.datab(data_out_11),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\max[11]~11_combout ),
	.cout());
defparam \max[11]~11 .lut_mask = 16'hAACC;
defparam \max[11]~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \max[11]~12 (
	.dataa(\Add0~22_combout ),
	.datab(\Add1~22_combout ),
	.datac(gnd),
	.datad(\LessThan0~22_combout ),
	.cin(gnd),
	.combout(\max[11]~12_combout ),
	.cout());
defparam \max[11]~12 .lut_mask = 16'hAACC;
defparam \max[11]~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mag_reg[11]~35 (
	.dataa(\max[11]~11_combout ),
	.datab(\max[11]~12_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\mag_reg[10]~34 ),
	.combout(\mag_reg[11]~35_combout ),
	.cout(\mag_reg[11]~36 ));
defparam \mag_reg[11]~35 .lut_mask = 16'h787F;
defparam \mag_reg[11]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \mag_reg[12]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\mag_reg[11]~36 ),
	.combout(\mag_reg[12]~37_combout ),
	.cout());
defparam \mag_reg[12]~37 .lut_mask = 16'h0F0F;
defparam \mag_reg[12]~37 .sum_lutc_input = "cin";

endmodule

module lms_dsp_counter (
	count_reg_0,
	running_reg1,
	count_reg_1,
	count_reg_2,
	count_reg_3,
	count_reg_4,
	count_reg_5,
	count_reg_6,
	count_reg_7,
	count_reg_8,
	count_reg_9,
	count_reg_10,
	count_reg_11,
	count_reg_12,
	count_reg_13,
	count_reg_14,
	count_reg_15,
	altera_reset_synchronizer_int_chain_out,
	launch,
	delay_reg_24_1,
	clock,
	ppd_cfg_passthrough_len_15,
	ppd_cfg_passthrough_len_14,
	ppd_cfg_passthrough_len_13,
	ppd_cfg_passthrough_len_12,
	ppd_cfg_passthrough_len_11,
	ppd_cfg_passthrough_len_10,
	ppd_cfg_passthrough_len_9,
	ppd_cfg_passthrough_len_8,
	ppd_cfg_passthrough_len_7,
	ppd_cfg_passthrough_len_6,
	ppd_cfg_passthrough_len_5,
	ppd_cfg_passthrough_len_4,
	ppd_cfg_passthrough_len_3,
	ppd_cfg_passthrough_len_2,
	ppd_cfg_passthrough_len_1,
	ppd_cfg_passthrough_len_0)/* synthesis synthesis_greybox=0 */;
output 	count_reg_0;
output 	running_reg1;
output 	count_reg_1;
output 	count_reg_2;
output 	count_reg_3;
output 	count_reg_4;
output 	count_reg_5;
output 	count_reg_6;
output 	count_reg_7;
output 	count_reg_8;
output 	count_reg_9;
output 	count_reg_10;
output 	count_reg_11;
output 	count_reg_12;
output 	count_reg_13;
output 	count_reg_14;
output 	count_reg_15;
input 	altera_reset_synchronizer_int_chain_out;
input 	launch;
input 	delay_reg_24_1;
input 	clock;
input 	ppd_cfg_passthrough_len_15;
input 	ppd_cfg_passthrough_len_14;
input 	ppd_cfg_passthrough_len_13;
input 	ppd_cfg_passthrough_len_12;
input 	ppd_cfg_passthrough_len_11;
input 	ppd_cfg_passthrough_len_10;
input 	ppd_cfg_passthrough_len_9;
input 	ppd_cfg_passthrough_len_8;
input 	ppd_cfg_passthrough_len_7;
input 	ppd_cfg_passthrough_len_6;
input 	ppd_cfg_passthrough_len_5;
input 	ppd_cfg_passthrough_len_4;
input 	ppd_cfg_passthrough_len_3;
input 	ppd_cfg_passthrough_len_2;
input 	ppd_cfg_passthrough_len_1;
input 	ppd_cfg_passthrough_len_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~0_combout ;
wire \LessThan1~1_cout ;
wire \LessThan1~3_cout ;
wire \LessThan1~5_cout ;
wire \LessThan1~7_cout ;
wire \LessThan1~9_cout ;
wire \LessThan1~11_cout ;
wire \LessThan1~13_cout ;
wire \LessThan1~15_cout ;
wire \LessThan1~17_cout ;
wire \LessThan1~19_cout ;
wire \LessThan1~21_cout ;
wire \LessThan1~23_cout ;
wire \LessThan1~25_cout ;
wire \LessThan1~27_cout ;
wire \LessThan1~29_cout ;
wire \LessThan1~30_combout ;
wire \always0~0_combout ;
wire \always0~1_combout ;
wire \always0~2_combout ;
wire \always0~3_combout ;
wire \always0~4_combout ;
wire \count_reg~0_combout ;
wire \running_reg~0_combout ;
wire \running_reg~1_combout ;
wire \count_reg[2]~1_combout ;
wire \Add0~1 ;
wire \Add0~2_combout ;
wire \count_reg~2_combout ;
wire \Add0~3 ;
wire \Add0~4_combout ;
wire \count_reg~3_combout ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \count_reg~4_combout ;
wire \Add0~7 ;
wire \Add0~8_combout ;
wire \count_reg~5_combout ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \count_reg~6_combout ;
wire \Add0~11 ;
wire \Add0~12_combout ;
wire \count_reg~7_combout ;
wire \Add0~13 ;
wire \Add0~14_combout ;
wire \count_reg~8_combout ;
wire \Add0~15 ;
wire \Add0~16_combout ;
wire \count_reg~9_combout ;
wire \Add0~17 ;
wire \Add0~18_combout ;
wire \count_reg~10_combout ;
wire \Add0~19 ;
wire \Add0~20_combout ;
wire \count_reg~11_combout ;
wire \Add0~21 ;
wire \Add0~22_combout ;
wire \count_reg~12_combout ;
wire \Add0~23 ;
wire \Add0~24_combout ;
wire \count_reg~13_combout ;
wire \Add0~25 ;
wire \Add0~26_combout ;
wire \count_reg~14_combout ;
wire \Add0~27 ;
wire \Add0~28_combout ;
wire \count_reg~15_combout ;
wire \Add0~29 ;
wire \Add0~30_combout ;
wire \count_reg~16_combout ;


dffeas \count_reg[0] (
	.clk(clock),
	.d(\count_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(\running_reg~0_combout ),
	.q(count_reg_0),
	.prn(vcc));
defparam \count_reg[0] .is_wysiwyg = "true";
defparam \count_reg[0] .power_up = "low";

dffeas running_reg(
	.clk(clock),
	.d(\running_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(\running_reg~0_combout ),
	.q(running_reg1),
	.prn(vcc));
defparam running_reg.is_wysiwyg = "true";
defparam running_reg.power_up = "low";

dffeas \count_reg[1] (
	.clk(clock),
	.d(\count_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\running_reg~0_combout ),
	.q(count_reg_1),
	.prn(vcc));
defparam \count_reg[1] .is_wysiwyg = "true";
defparam \count_reg[1] .power_up = "low";

dffeas \count_reg[2] (
	.clk(clock),
	.d(\count_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\running_reg~0_combout ),
	.q(count_reg_2),
	.prn(vcc));
defparam \count_reg[2] .is_wysiwyg = "true";
defparam \count_reg[2] .power_up = "low";

dffeas \count_reg[3] (
	.clk(clock),
	.d(\count_reg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\running_reg~0_combout ),
	.q(count_reg_3),
	.prn(vcc));
defparam \count_reg[3] .is_wysiwyg = "true";
defparam \count_reg[3] .power_up = "low";

dffeas \count_reg[4] (
	.clk(clock),
	.d(\count_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\running_reg~0_combout ),
	.q(count_reg_4),
	.prn(vcc));
defparam \count_reg[4] .is_wysiwyg = "true";
defparam \count_reg[4] .power_up = "low";

dffeas \count_reg[5] (
	.clk(clock),
	.d(\count_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\running_reg~0_combout ),
	.q(count_reg_5),
	.prn(vcc));
defparam \count_reg[5] .is_wysiwyg = "true";
defparam \count_reg[5] .power_up = "low";

dffeas \count_reg[6] (
	.clk(clock),
	.d(\count_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\running_reg~0_combout ),
	.q(count_reg_6),
	.prn(vcc));
defparam \count_reg[6] .is_wysiwyg = "true";
defparam \count_reg[6] .power_up = "low";

dffeas \count_reg[7] (
	.clk(clock),
	.d(\count_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\running_reg~0_combout ),
	.q(count_reg_7),
	.prn(vcc));
defparam \count_reg[7] .is_wysiwyg = "true";
defparam \count_reg[7] .power_up = "low";

dffeas \count_reg[8] (
	.clk(clock),
	.d(\count_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\running_reg~0_combout ),
	.q(count_reg_8),
	.prn(vcc));
defparam \count_reg[8] .is_wysiwyg = "true";
defparam \count_reg[8] .power_up = "low";

dffeas \count_reg[9] (
	.clk(clock),
	.d(\count_reg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\running_reg~0_combout ),
	.q(count_reg_9),
	.prn(vcc));
defparam \count_reg[9] .is_wysiwyg = "true";
defparam \count_reg[9] .power_up = "low";

dffeas \count_reg[10] (
	.clk(clock),
	.d(\count_reg~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\running_reg~0_combout ),
	.q(count_reg_10),
	.prn(vcc));
defparam \count_reg[10] .is_wysiwyg = "true";
defparam \count_reg[10] .power_up = "low";

dffeas \count_reg[11] (
	.clk(clock),
	.d(\count_reg~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\running_reg~0_combout ),
	.q(count_reg_11),
	.prn(vcc));
defparam \count_reg[11] .is_wysiwyg = "true";
defparam \count_reg[11] .power_up = "low";

dffeas \count_reg[12] (
	.clk(clock),
	.d(\count_reg~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\running_reg~0_combout ),
	.q(count_reg_12),
	.prn(vcc));
defparam \count_reg[12] .is_wysiwyg = "true";
defparam \count_reg[12] .power_up = "low";

dffeas \count_reg[13] (
	.clk(clock),
	.d(\count_reg~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\running_reg~0_combout ),
	.q(count_reg_13),
	.prn(vcc));
defparam \count_reg[13] .is_wysiwyg = "true";
defparam \count_reg[13] .power_up = "low";

dffeas \count_reg[14] (
	.clk(clock),
	.d(\count_reg~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\running_reg~0_combout ),
	.q(count_reg_14),
	.prn(vcc));
defparam \count_reg[14] .is_wysiwyg = "true";
defparam \count_reg[14] .power_up = "low";

dffeas \count_reg[15] (
	.clk(clock),
	.d(\count_reg~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\running_reg~0_combout ),
	.q(count_reg_15),
	.prn(vcc));
defparam \count_reg[15] .is_wysiwyg = "true";
defparam \count_reg[15] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~0 (
	.dataa(count_reg_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
defparam \Add0~0 .lut_mask = 16'h55AA;
defparam \Add0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \LessThan1~1 (
	.dataa(count_reg_0),
	.datab(ppd_cfg_passthrough_len_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan1~1_cout ));
defparam \LessThan1~1 .lut_mask = 16'h0044;
defparam \LessThan1~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan1~3 (
	.dataa(count_reg_1),
	.datab(ppd_cfg_passthrough_len_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~1_cout ),
	.combout(),
	.cout(\LessThan1~3_cout ));
defparam \LessThan1~3 .lut_mask = 16'h002B;
defparam \LessThan1~3 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan1~5 (
	.dataa(count_reg_2),
	.datab(ppd_cfg_passthrough_len_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~3_cout ),
	.combout(),
	.cout(\LessThan1~5_cout ));
defparam \LessThan1~5 .lut_mask = 16'h004D;
defparam \LessThan1~5 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan1~7 (
	.dataa(count_reg_3),
	.datab(ppd_cfg_passthrough_len_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~5_cout ),
	.combout(),
	.cout(\LessThan1~7_cout ));
defparam \LessThan1~7 .lut_mask = 16'h002B;
defparam \LessThan1~7 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan1~9 (
	.dataa(count_reg_4),
	.datab(ppd_cfg_passthrough_len_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~7_cout ),
	.combout(),
	.cout(\LessThan1~9_cout ));
defparam \LessThan1~9 .lut_mask = 16'h004D;
defparam \LessThan1~9 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan1~11 (
	.dataa(count_reg_5),
	.datab(ppd_cfg_passthrough_len_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~9_cout ),
	.combout(),
	.cout(\LessThan1~11_cout ));
defparam \LessThan1~11 .lut_mask = 16'h002B;
defparam \LessThan1~11 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan1~13 (
	.dataa(count_reg_6),
	.datab(ppd_cfg_passthrough_len_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~11_cout ),
	.combout(),
	.cout(\LessThan1~13_cout ));
defparam \LessThan1~13 .lut_mask = 16'h004D;
defparam \LessThan1~13 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan1~15 (
	.dataa(count_reg_7),
	.datab(ppd_cfg_passthrough_len_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~13_cout ),
	.combout(),
	.cout(\LessThan1~15_cout ));
defparam \LessThan1~15 .lut_mask = 16'h002B;
defparam \LessThan1~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan1~17 (
	.dataa(count_reg_8),
	.datab(ppd_cfg_passthrough_len_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~15_cout ),
	.combout(),
	.cout(\LessThan1~17_cout ));
defparam \LessThan1~17 .lut_mask = 16'h004D;
defparam \LessThan1~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan1~19 (
	.dataa(count_reg_9),
	.datab(ppd_cfg_passthrough_len_9),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~17_cout ),
	.combout(),
	.cout(\LessThan1~19_cout ));
defparam \LessThan1~19 .lut_mask = 16'h002B;
defparam \LessThan1~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan1~21 (
	.dataa(count_reg_10),
	.datab(ppd_cfg_passthrough_len_10),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~19_cout ),
	.combout(),
	.cout(\LessThan1~21_cout ));
defparam \LessThan1~21 .lut_mask = 16'h004D;
defparam \LessThan1~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan1~23 (
	.dataa(count_reg_11),
	.datab(ppd_cfg_passthrough_len_11),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~21_cout ),
	.combout(),
	.cout(\LessThan1~23_cout ));
defparam \LessThan1~23 .lut_mask = 16'h002B;
defparam \LessThan1~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan1~25 (
	.dataa(count_reg_12),
	.datab(ppd_cfg_passthrough_len_12),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~23_cout ),
	.combout(),
	.cout(\LessThan1~25_cout ));
defparam \LessThan1~25 .lut_mask = 16'h004D;
defparam \LessThan1~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan1~27 (
	.dataa(count_reg_13),
	.datab(ppd_cfg_passthrough_len_13),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~25_cout ),
	.combout(),
	.cout(\LessThan1~27_cout ));
defparam \LessThan1~27 .lut_mask = 16'h002B;
defparam \LessThan1~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan1~29 (
	.dataa(count_reg_14),
	.datab(ppd_cfg_passthrough_len_14),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~27_cout ),
	.combout(),
	.cout(\LessThan1~29_cout ));
defparam \LessThan1~29 .lut_mask = 16'h004D;
defparam \LessThan1~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan1~30 (
	.dataa(count_reg_15),
	.datab(ppd_cfg_passthrough_len_15),
	.datac(gnd),
	.datad(gnd),
	.cin(\LessThan1~29_cout ),
	.combout(\LessThan1~30_combout ),
	.cout());
defparam \LessThan1~30 .lut_mask = 16'hD4D4;
defparam \LessThan1~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \always0~0 (
	.dataa(count_reg_1),
	.datab(count_reg_2),
	.datac(count_reg_3),
	.datad(count_reg_4),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'h0001;
defparam \always0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always0~1 (
	.dataa(count_reg_5),
	.datab(count_reg_6),
	.datac(count_reg_7),
	.datad(count_reg_8),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
defparam \always0~1 .lut_mask = 16'h0001;
defparam \always0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always0~2 (
	.dataa(count_reg_9),
	.datab(count_reg_10),
	.datac(count_reg_11),
	.datad(count_reg_12),
	.cin(gnd),
	.combout(\always0~2_combout ),
	.cout());
defparam \always0~2 .lut_mask = 16'h0001;
defparam \always0~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always0~3 (
	.dataa(count_reg_0),
	.datab(count_reg_13),
	.datac(count_reg_14),
	.datad(count_reg_15),
	.cin(gnd),
	.combout(\always0~3_combout ),
	.cout());
defparam \always0~3 .lut_mask = 16'h0001;
defparam \always0~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always0~4 (
	.dataa(\always0~0_combout ),
	.datab(\always0~1_combout ),
	.datac(\always0~2_combout ),
	.datad(\always0~3_combout ),
	.cin(gnd),
	.combout(\always0~4_combout ),
	.cout());
defparam \always0~4 .lut_mask = 16'h8000;
defparam \always0~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \count_reg~0 (
	.dataa(\Add0~0_combout ),
	.datab(launch),
	.datac(\LessThan1~30_combout ),
	.datad(\always0~4_combout ),
	.cin(gnd),
	.combout(\count_reg~0_combout ),
	.cout());
defparam \count_reg~0 .lut_mask = 16'h88AC;
defparam \count_reg~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \running_reg~0 (
	.dataa(delay_reg_24_1),
	.datab(gnd),
	.datac(gnd),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\running_reg~0_combout ),
	.cout());
defparam \running_reg~0 .lut_mask = 16'hAAFF;
defparam \running_reg~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \running_reg~1 (
	.dataa(launch),
	.datab(\LessThan1~30_combout ),
	.datac(gnd),
	.datad(\always0~4_combout ),
	.cin(gnd),
	.combout(\running_reg~1_combout ),
	.cout());
defparam \running_reg~1 .lut_mask = 16'hAAEE;
defparam \running_reg~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \count_reg[2]~1 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(launch),
	.datac(\LessThan1~30_combout ),
	.datad(\always0~4_combout ),
	.cin(gnd),
	.combout(\count_reg[2]~1_combout ),
	.cout());
defparam \count_reg[2]~1 .lut_mask = 16'h88A0;
defparam \count_reg[2]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~2 (
	.dataa(count_reg_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'h5A5F;
defparam \Add0~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count_reg~2 (
	.dataa(\count_reg[2]~1_combout ),
	.datab(\Add0~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count_reg~2_combout ),
	.cout());
defparam \count_reg~2 .lut_mask = 16'h8888;
defparam \count_reg~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~4 (
	.dataa(count_reg_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'hA50A;
defparam \Add0~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count_reg~3 (
	.dataa(\count_reg[2]~1_combout ),
	.datab(\Add0~4_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count_reg~3_combout ),
	.cout());
defparam \count_reg~3 .lut_mask = 16'h8888;
defparam \count_reg~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~6 (
	.dataa(count_reg_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'h5A5F;
defparam \Add0~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count_reg~4 (
	.dataa(\count_reg[2]~1_combout ),
	.datab(\Add0~6_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count_reg~4_combout ),
	.cout());
defparam \count_reg~4 .lut_mask = 16'h8888;
defparam \count_reg~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~8 (
	.dataa(count_reg_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
defparam \Add0~8 .lut_mask = 16'hA50A;
defparam \Add0~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count_reg~5 (
	.dataa(\count_reg[2]~1_combout ),
	.datab(\Add0~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count_reg~5_combout ),
	.cout());
defparam \count_reg~5 .lut_mask = 16'h8888;
defparam \count_reg~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~10 (
	.dataa(count_reg_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
defparam \Add0~10 .lut_mask = 16'h5A5F;
defparam \Add0~10 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count_reg~6 (
	.dataa(\count_reg[2]~1_combout ),
	.datab(\Add0~10_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count_reg~6_combout ),
	.cout());
defparam \count_reg~6 .lut_mask = 16'h8888;
defparam \count_reg~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~12 (
	.dataa(count_reg_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
defparam \Add0~12 .lut_mask = 16'hA50A;
defparam \Add0~12 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count_reg~7 (
	.dataa(\count_reg[2]~1_combout ),
	.datab(\Add0~12_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count_reg~7_combout ),
	.cout());
defparam \count_reg~7 .lut_mask = 16'h8888;
defparam \count_reg~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~14 (
	.dataa(count_reg_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
defparam \Add0~14 .lut_mask = 16'h5A5F;
defparam \Add0~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count_reg~8 (
	.dataa(\count_reg[2]~1_combout ),
	.datab(\Add0~14_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count_reg~8_combout ),
	.cout());
defparam \count_reg~8 .lut_mask = 16'h8888;
defparam \count_reg~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~16 (
	.dataa(count_reg_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout(\Add0~17 ));
defparam \Add0~16 .lut_mask = 16'hA50A;
defparam \Add0~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count_reg~9 (
	.dataa(\count_reg[2]~1_combout ),
	.datab(\Add0~16_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count_reg~9_combout ),
	.cout());
defparam \count_reg~9 .lut_mask = 16'h8888;
defparam \count_reg~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~18 (
	.dataa(count_reg_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~17 ),
	.combout(\Add0~18_combout ),
	.cout(\Add0~19 ));
defparam \Add0~18 .lut_mask = 16'h5A5F;
defparam \Add0~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count_reg~10 (
	.dataa(\count_reg[2]~1_combout ),
	.datab(\Add0~18_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count_reg~10_combout ),
	.cout());
defparam \count_reg~10 .lut_mask = 16'h8888;
defparam \count_reg~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~20 (
	.dataa(count_reg_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~19 ),
	.combout(\Add0~20_combout ),
	.cout(\Add0~21 ));
defparam \Add0~20 .lut_mask = 16'hA50A;
defparam \Add0~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count_reg~11 (
	.dataa(\count_reg[2]~1_combout ),
	.datab(\Add0~20_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count_reg~11_combout ),
	.cout());
defparam \count_reg~11 .lut_mask = 16'h8888;
defparam \count_reg~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~22 (
	.dataa(count_reg_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~21 ),
	.combout(\Add0~22_combout ),
	.cout(\Add0~23 ));
defparam \Add0~22 .lut_mask = 16'h5A5F;
defparam \Add0~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count_reg~12 (
	.dataa(\count_reg[2]~1_combout ),
	.datab(\Add0~22_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count_reg~12_combout ),
	.cout());
defparam \count_reg~12 .lut_mask = 16'h8888;
defparam \count_reg~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~24 (
	.dataa(count_reg_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~23 ),
	.combout(\Add0~24_combout ),
	.cout(\Add0~25 ));
defparam \Add0~24 .lut_mask = 16'hA50A;
defparam \Add0~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count_reg~13 (
	.dataa(\count_reg[2]~1_combout ),
	.datab(\Add0~24_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count_reg~13_combout ),
	.cout());
defparam \count_reg~13 .lut_mask = 16'h8888;
defparam \count_reg~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~26 (
	.dataa(count_reg_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~25 ),
	.combout(\Add0~26_combout ),
	.cout(\Add0~27 ));
defparam \Add0~26 .lut_mask = 16'h5A5F;
defparam \Add0~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count_reg~14 (
	.dataa(\count_reg[2]~1_combout ),
	.datab(\Add0~26_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count_reg~14_combout ),
	.cout());
defparam \count_reg~14 .lut_mask = 16'h8888;
defparam \count_reg~14 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~28 (
	.dataa(count_reg_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~27 ),
	.combout(\Add0~28_combout ),
	.cout(\Add0~29 ));
defparam \Add0~28 .lut_mask = 16'hA50A;
defparam \Add0~28 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count_reg~15 (
	.dataa(\count_reg[2]~1_combout ),
	.datab(\Add0~28_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count_reg~15_combout ),
	.cout());
defparam \count_reg~15 .lut_mask = 16'h8888;
defparam \count_reg~15 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~30 (
	.dataa(count_reg_15),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~29 ),
	.combout(\Add0~30_combout ),
	.cout());
defparam \Add0~30 .lut_mask = 16'h5A5A;
defparam \Add0~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count_reg~16 (
	.dataa(\count_reg[2]~1_combout ),
	.datab(\Add0~30_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count_reg~16_combout ),
	.cout());
defparam \count_reg~16 .lut_mask = 16'h8888;
defparam \count_reg~16 .sum_lutc_input = "datac";

endmodule

module lms_dsp_delay_line (
	altera_reset_synchronizer_int_chain_out,
	delay_reg_24_1,
	delay_reg_24_0,
	data_out_12,
	data_out_0,
	data_out_11,
	data_out_10,
	data_out_9,
	data_out_8,
	data_out_7,
	data_out_6,
	data_out_5,
	data_out_4,
	data_out_3,
	data_out_2,
	data_out_1,
	data_out_23,
	data_out_22,
	data_out_21,
	data_out_20,
	data_out_19,
	data_out_18,
	data_out_17,
	data_out_16,
	data_out_15,
	data_out_14,
	data_out_13,
	data_valid,
	delay_reg_25_2,
	delay_reg_0_3,
	delay_reg_1_3,
	delay_reg_2_3,
	delay_reg_3_3,
	delay_reg_4_3,
	delay_reg_5_3,
	delay_reg_6_3,
	delay_reg_7_3,
	delay_reg_8_3,
	delay_reg_9_3,
	delay_reg_10_3,
	delay_reg_11_3,
	delay_reg_12_3,
	delay_reg_13_3,
	delay_reg_14_3,
	delay_reg_15_3,
	delay_reg_16_3,
	delay_reg_17_3,
	delay_reg_18_3,
	delay_reg_19_3,
	delay_reg_20_3,
	delay_reg_21_3,
	delay_reg_22_3,
	delay_reg_23_3,
	delay_reg_24_3,
	clock,
	ppd_cfg_enable)/* synthesis synthesis_greybox=0 */;
input 	altera_reset_synchronizer_int_chain_out;
output 	delay_reg_24_1;
output 	delay_reg_24_0;
input 	data_out_12;
input 	data_out_0;
input 	data_out_11;
input 	data_out_10;
input 	data_out_9;
input 	data_out_8;
input 	data_out_7;
input 	data_out_6;
input 	data_out_5;
input 	data_out_4;
input 	data_out_3;
input 	data_out_2;
input 	data_out_1;
input 	data_out_23;
input 	data_out_22;
input 	data_out_21;
input 	data_out_20;
input 	data_out_19;
input 	data_out_18;
input 	data_out_17;
input 	data_out_16;
input 	data_out_15;
input 	data_out_14;
input 	data_out_13;
input 	data_valid;
output 	delay_reg_25_2;
output 	delay_reg_0_3;
output 	delay_reg_1_3;
output 	delay_reg_2_3;
output 	delay_reg_3_3;
output 	delay_reg_4_3;
output 	delay_reg_5_3;
output 	delay_reg_6_3;
output 	delay_reg_7_3;
output 	delay_reg_8_3;
output 	delay_reg_9_3;
output 	delay_reg_10_3;
output 	delay_reg_11_3;
output 	delay_reg_12_3;
output 	delay_reg_13_3;
output 	delay_reg_14_3;
output 	delay_reg_15_3;
output 	delay_reg_16_3;
output 	delay_reg_17_3;
output 	delay_reg_18_3;
output 	delay_reg_19_3;
output 	delay_reg_20_3;
output 	delay_reg_21_3;
output 	delay_reg_22_3;
output 	delay_reg_23_3;
output 	delay_reg_24_3;
input 	clock;
input 	ppd_cfg_enable;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \delay_reg~0_combout ;
wire \delay_reg~1_combout ;
wire \delay_reg~54_combout ;
wire \delay_reg[0][25]~q ;
wire \delay_reg~28_combout ;
wire \delay_reg[1][25]~q ;
wire \delay_reg~2_combout ;
wire \delay_reg~79_combout ;
wire \delay_reg[0][0]~q ;
wire \delay_reg~55_combout ;
wire \delay_reg[1][0]~q ;
wire \delay_reg~29_combout ;
wire \delay_reg[2][0]~q ;
wire \delay_reg~3_combout ;
wire \delay_reg~80_combout ;
wire \delay_reg[0][1]~q ;
wire \delay_reg~56_combout ;
wire \delay_reg[1][1]~q ;
wire \delay_reg~30_combout ;
wire \delay_reg[2][1]~q ;
wire \delay_reg~4_combout ;
wire \delay_reg~81_combout ;
wire \delay_reg[0][2]~q ;
wire \delay_reg~57_combout ;
wire \delay_reg[1][2]~q ;
wire \delay_reg~31_combout ;
wire \delay_reg[2][2]~q ;
wire \delay_reg~5_combout ;
wire \delay_reg~82_combout ;
wire \delay_reg[0][3]~q ;
wire \delay_reg~58_combout ;
wire \delay_reg[1][3]~q ;
wire \delay_reg~32_combout ;
wire \delay_reg[2][3]~q ;
wire \delay_reg~6_combout ;
wire \delay_reg~83_combout ;
wire \delay_reg[0][4]~q ;
wire \delay_reg~59_combout ;
wire \delay_reg[1][4]~q ;
wire \delay_reg~33_combout ;
wire \delay_reg[2][4]~q ;
wire \delay_reg~7_combout ;
wire \delay_reg~84_combout ;
wire \delay_reg[0][5]~q ;
wire \delay_reg~60_combout ;
wire \delay_reg[1][5]~q ;
wire \delay_reg~34_combout ;
wire \delay_reg[2][5]~q ;
wire \delay_reg~8_combout ;
wire \delay_reg~85_combout ;
wire \delay_reg[0][6]~q ;
wire \delay_reg~61_combout ;
wire \delay_reg[1][6]~q ;
wire \delay_reg~35_combout ;
wire \delay_reg[2][6]~q ;
wire \delay_reg~9_combout ;
wire \delay_reg~86_combout ;
wire \delay_reg[0][7]~q ;
wire \delay_reg~62_combout ;
wire \delay_reg[1][7]~q ;
wire \delay_reg~36_combout ;
wire \delay_reg[2][7]~q ;
wire \delay_reg~10_combout ;
wire \delay_reg~87_combout ;
wire \delay_reg[0][8]~q ;
wire \delay_reg~63_combout ;
wire \delay_reg[1][8]~q ;
wire \delay_reg~37_combout ;
wire \delay_reg[2][8]~q ;
wire \delay_reg~11_combout ;
wire \delay_reg~88_combout ;
wire \delay_reg[0][9]~q ;
wire \delay_reg~64_combout ;
wire \delay_reg[1][9]~q ;
wire \delay_reg~38_combout ;
wire \delay_reg[2][9]~q ;
wire \delay_reg~12_combout ;
wire \delay_reg~89_combout ;
wire \delay_reg[0][10]~q ;
wire \delay_reg~65_combout ;
wire \delay_reg[1][10]~q ;
wire \delay_reg~39_combout ;
wire \delay_reg[2][10]~q ;
wire \delay_reg~13_combout ;
wire \delay_reg~90_combout ;
wire \delay_reg[0][11]~q ;
wire \delay_reg~66_combout ;
wire \delay_reg[1][11]~q ;
wire \delay_reg~40_combout ;
wire \delay_reg[2][11]~q ;
wire \delay_reg~14_combout ;
wire \delay_reg~91_combout ;
wire \delay_reg[0][12]~q ;
wire \delay_reg~67_combout ;
wire \delay_reg[1][12]~q ;
wire \delay_reg~41_combout ;
wire \delay_reg[2][12]~q ;
wire \delay_reg~15_combout ;
wire \delay_reg~92_combout ;
wire \delay_reg[0][13]~q ;
wire \delay_reg~68_combout ;
wire \delay_reg[1][13]~q ;
wire \delay_reg~42_combout ;
wire \delay_reg[2][13]~q ;
wire \delay_reg~16_combout ;
wire \delay_reg~93_combout ;
wire \delay_reg[0][14]~q ;
wire \delay_reg~69_combout ;
wire \delay_reg[1][14]~q ;
wire \delay_reg~43_combout ;
wire \delay_reg[2][14]~q ;
wire \delay_reg~17_combout ;
wire \delay_reg~94_combout ;
wire \delay_reg[0][15]~q ;
wire \delay_reg~70_combout ;
wire \delay_reg[1][15]~q ;
wire \delay_reg~44_combout ;
wire \delay_reg[2][15]~q ;
wire \delay_reg~18_combout ;
wire \delay_reg~95_combout ;
wire \delay_reg[0][16]~q ;
wire \delay_reg~71_combout ;
wire \delay_reg[1][16]~q ;
wire \delay_reg~45_combout ;
wire \delay_reg[2][16]~q ;
wire \delay_reg~19_combout ;
wire \delay_reg~96_combout ;
wire \delay_reg[0][17]~q ;
wire \delay_reg~72_combout ;
wire \delay_reg[1][17]~q ;
wire \delay_reg~46_combout ;
wire \delay_reg[2][17]~q ;
wire \delay_reg~20_combout ;
wire \delay_reg~97_combout ;
wire \delay_reg[0][18]~q ;
wire \delay_reg~73_combout ;
wire \delay_reg[1][18]~q ;
wire \delay_reg~47_combout ;
wire \delay_reg[2][18]~q ;
wire \delay_reg~21_combout ;
wire \delay_reg~98_combout ;
wire \delay_reg[0][19]~q ;
wire \delay_reg~74_combout ;
wire \delay_reg[1][19]~q ;
wire \delay_reg~48_combout ;
wire \delay_reg[2][19]~q ;
wire \delay_reg~22_combout ;
wire \delay_reg~99_combout ;
wire \delay_reg[0][20]~q ;
wire \delay_reg~75_combout ;
wire \delay_reg[1][20]~q ;
wire \delay_reg~49_combout ;
wire \delay_reg[2][20]~q ;
wire \delay_reg~23_combout ;
wire \delay_reg~100_combout ;
wire \delay_reg[0][21]~q ;
wire \delay_reg~76_combout ;
wire \delay_reg[1][21]~q ;
wire \delay_reg~50_combout ;
wire \delay_reg[2][21]~q ;
wire \delay_reg~24_combout ;
wire \delay_reg~101_combout ;
wire \delay_reg[0][22]~q ;
wire \delay_reg~77_combout ;
wire \delay_reg[1][22]~q ;
wire \delay_reg~51_combout ;
wire \delay_reg[2][22]~q ;
wire \delay_reg~25_combout ;
wire \delay_reg~102_combout ;
wire \delay_reg[0][23]~q ;
wire \delay_reg~78_combout ;
wire \delay_reg[1][23]~q ;
wire \delay_reg~52_combout ;
wire \delay_reg[2][23]~q ;
wire \delay_reg~26_combout ;
wire \delay_reg~53_combout ;
wire \delay_reg[2][24]~q ;
wire \delay_reg~27_combout ;


dffeas \delay_reg[1][24] (
	.clk(clock),
	.d(\delay_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_24_1),
	.prn(vcc));
defparam \delay_reg[1][24] .is_wysiwyg = "true";
defparam \delay_reg[1][24] .power_up = "low";

dffeas \delay_reg[0][24] (
	.clk(clock),
	.d(\delay_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_24_0),
	.prn(vcc));
defparam \delay_reg[0][24] .is_wysiwyg = "true";
defparam \delay_reg[0][24] .power_up = "low";

dffeas \delay_reg[2][25] (
	.clk(clock),
	.d(\delay_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_25_2),
	.prn(vcc));
defparam \delay_reg[2][25] .is_wysiwyg = "true";
defparam \delay_reg[2][25] .power_up = "low";

dffeas \delay_reg[3][0] (
	.clk(clock),
	.d(\delay_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_0_3),
	.prn(vcc));
defparam \delay_reg[3][0] .is_wysiwyg = "true";
defparam \delay_reg[3][0] .power_up = "low";

dffeas \delay_reg[3][1] (
	.clk(clock),
	.d(\delay_reg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_1_3),
	.prn(vcc));
defparam \delay_reg[3][1] .is_wysiwyg = "true";
defparam \delay_reg[3][1] .power_up = "low";

dffeas \delay_reg[3][2] (
	.clk(clock),
	.d(\delay_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_2_3),
	.prn(vcc));
defparam \delay_reg[3][2] .is_wysiwyg = "true";
defparam \delay_reg[3][2] .power_up = "low";

dffeas \delay_reg[3][3] (
	.clk(clock),
	.d(\delay_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_3_3),
	.prn(vcc));
defparam \delay_reg[3][3] .is_wysiwyg = "true";
defparam \delay_reg[3][3] .power_up = "low";

dffeas \delay_reg[3][4] (
	.clk(clock),
	.d(\delay_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_4_3),
	.prn(vcc));
defparam \delay_reg[3][4] .is_wysiwyg = "true";
defparam \delay_reg[3][4] .power_up = "low";

dffeas \delay_reg[3][5] (
	.clk(clock),
	.d(\delay_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_5_3),
	.prn(vcc));
defparam \delay_reg[3][5] .is_wysiwyg = "true";
defparam \delay_reg[3][5] .power_up = "low";

dffeas \delay_reg[3][6] (
	.clk(clock),
	.d(\delay_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_6_3),
	.prn(vcc));
defparam \delay_reg[3][6] .is_wysiwyg = "true";
defparam \delay_reg[3][6] .power_up = "low";

dffeas \delay_reg[3][7] (
	.clk(clock),
	.d(\delay_reg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_7_3),
	.prn(vcc));
defparam \delay_reg[3][7] .is_wysiwyg = "true";
defparam \delay_reg[3][7] .power_up = "low";

dffeas \delay_reg[3][8] (
	.clk(clock),
	.d(\delay_reg~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_8_3),
	.prn(vcc));
defparam \delay_reg[3][8] .is_wysiwyg = "true";
defparam \delay_reg[3][8] .power_up = "low";

dffeas \delay_reg[3][9] (
	.clk(clock),
	.d(\delay_reg~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_9_3),
	.prn(vcc));
defparam \delay_reg[3][9] .is_wysiwyg = "true";
defparam \delay_reg[3][9] .power_up = "low";

dffeas \delay_reg[3][10] (
	.clk(clock),
	.d(\delay_reg~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_10_3),
	.prn(vcc));
defparam \delay_reg[3][10] .is_wysiwyg = "true";
defparam \delay_reg[3][10] .power_up = "low";

dffeas \delay_reg[3][11] (
	.clk(clock),
	.d(\delay_reg~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_11_3),
	.prn(vcc));
defparam \delay_reg[3][11] .is_wysiwyg = "true";
defparam \delay_reg[3][11] .power_up = "low";

dffeas \delay_reg[3][12] (
	.clk(clock),
	.d(\delay_reg~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_12_3),
	.prn(vcc));
defparam \delay_reg[3][12] .is_wysiwyg = "true";
defparam \delay_reg[3][12] .power_up = "low";

dffeas \delay_reg[3][13] (
	.clk(clock),
	.d(\delay_reg~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_13_3),
	.prn(vcc));
defparam \delay_reg[3][13] .is_wysiwyg = "true";
defparam \delay_reg[3][13] .power_up = "low";

dffeas \delay_reg[3][14] (
	.clk(clock),
	.d(\delay_reg~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_14_3),
	.prn(vcc));
defparam \delay_reg[3][14] .is_wysiwyg = "true";
defparam \delay_reg[3][14] .power_up = "low";

dffeas \delay_reg[3][15] (
	.clk(clock),
	.d(\delay_reg~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_15_3),
	.prn(vcc));
defparam \delay_reg[3][15] .is_wysiwyg = "true";
defparam \delay_reg[3][15] .power_up = "low";

dffeas \delay_reg[3][16] (
	.clk(clock),
	.d(\delay_reg~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_16_3),
	.prn(vcc));
defparam \delay_reg[3][16] .is_wysiwyg = "true";
defparam \delay_reg[3][16] .power_up = "low";

dffeas \delay_reg[3][17] (
	.clk(clock),
	.d(\delay_reg~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_17_3),
	.prn(vcc));
defparam \delay_reg[3][17] .is_wysiwyg = "true";
defparam \delay_reg[3][17] .power_up = "low";

dffeas \delay_reg[3][18] (
	.clk(clock),
	.d(\delay_reg~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_18_3),
	.prn(vcc));
defparam \delay_reg[3][18] .is_wysiwyg = "true";
defparam \delay_reg[3][18] .power_up = "low";

dffeas \delay_reg[3][19] (
	.clk(clock),
	.d(\delay_reg~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_19_3),
	.prn(vcc));
defparam \delay_reg[3][19] .is_wysiwyg = "true";
defparam \delay_reg[3][19] .power_up = "low";

dffeas \delay_reg[3][20] (
	.clk(clock),
	.d(\delay_reg~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_20_3),
	.prn(vcc));
defparam \delay_reg[3][20] .is_wysiwyg = "true";
defparam \delay_reg[3][20] .power_up = "low";

dffeas \delay_reg[3][21] (
	.clk(clock),
	.d(\delay_reg~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_21_3),
	.prn(vcc));
defparam \delay_reg[3][21] .is_wysiwyg = "true";
defparam \delay_reg[3][21] .power_up = "low";

dffeas \delay_reg[3][22] (
	.clk(clock),
	.d(\delay_reg~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_22_3),
	.prn(vcc));
defparam \delay_reg[3][22] .is_wysiwyg = "true";
defparam \delay_reg[3][22] .power_up = "low";

dffeas \delay_reg[3][23] (
	.clk(clock),
	.d(\delay_reg~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_23_3),
	.prn(vcc));
defparam \delay_reg[3][23] .is_wysiwyg = "true";
defparam \delay_reg[3][23] .power_up = "low";

dffeas \delay_reg[3][24] (
	.clk(clock),
	.d(\delay_reg~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(delay_reg_24_3),
	.prn(vcc));
defparam \delay_reg[3][24] .is_wysiwyg = "true";
defparam \delay_reg[3][24] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(delay_reg_24_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~0_combout ),
	.cout());
defparam \delay_reg~0 .lut_mask = 16'h8888;
defparam \delay_reg~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~1 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_valid),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~1_combout ),
	.cout());
defparam \delay_reg~1 .lut_mask = 16'h8888;
defparam \delay_reg~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~54 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(ppd_cfg_enable),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~54_combout ),
	.cout());
defparam \delay_reg~54 .lut_mask = 16'h8888;
defparam \delay_reg~54 .sum_lutc_input = "datac";

dffeas \delay_reg[0][25] (
	.clk(clock),
	.d(\delay_reg~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][25]~q ),
	.prn(vcc));
defparam \delay_reg[0][25] .is_wysiwyg = "true";
defparam \delay_reg[0][25] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~28 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][25]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~28_combout ),
	.cout());
defparam \delay_reg~28 .lut_mask = 16'h8888;
defparam \delay_reg~28 .sum_lutc_input = "datac";

dffeas \delay_reg[1][25] (
	.clk(clock),
	.d(\delay_reg~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][25]~q ),
	.prn(vcc));
defparam \delay_reg[1][25] .is_wysiwyg = "true";
defparam \delay_reg[1][25] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~2 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][25]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~2_combout ),
	.cout());
defparam \delay_reg~2 .lut_mask = 16'h8888;
defparam \delay_reg~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~79 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~79_combout ),
	.cout());
defparam \delay_reg~79 .lut_mask = 16'h8888;
defparam \delay_reg~79 .sum_lutc_input = "datac";

dffeas \delay_reg[0][0] (
	.clk(clock),
	.d(\delay_reg~79_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][0]~q ),
	.prn(vcc));
defparam \delay_reg[0][0] .is_wysiwyg = "true";
defparam \delay_reg[0][0] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~55 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~55_combout ),
	.cout());
defparam \delay_reg~55 .lut_mask = 16'h8888;
defparam \delay_reg~55 .sum_lutc_input = "datac";

dffeas \delay_reg[1][0] (
	.clk(clock),
	.d(\delay_reg~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][0]~q ),
	.prn(vcc));
defparam \delay_reg[1][0] .is_wysiwyg = "true";
defparam \delay_reg[1][0] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~29 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~29_combout ),
	.cout());
defparam \delay_reg~29 .lut_mask = 16'h8888;
defparam \delay_reg~29 .sum_lutc_input = "datac";

dffeas \delay_reg[2][0] (
	.clk(clock),
	.d(\delay_reg~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][0]~q ),
	.prn(vcc));
defparam \delay_reg[2][0] .is_wysiwyg = "true";
defparam \delay_reg[2][0] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~3 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~3_combout ),
	.cout());
defparam \delay_reg~3 .lut_mask = 16'h8888;
defparam \delay_reg~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~80 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~80_combout ),
	.cout());
defparam \delay_reg~80 .lut_mask = 16'h8888;
defparam \delay_reg~80 .sum_lutc_input = "datac";

dffeas \delay_reg[0][1] (
	.clk(clock),
	.d(\delay_reg~80_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][1]~q ),
	.prn(vcc));
defparam \delay_reg[0][1] .is_wysiwyg = "true";
defparam \delay_reg[0][1] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~56 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~56_combout ),
	.cout());
defparam \delay_reg~56 .lut_mask = 16'h8888;
defparam \delay_reg~56 .sum_lutc_input = "datac";

dffeas \delay_reg[1][1] (
	.clk(clock),
	.d(\delay_reg~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][1]~q ),
	.prn(vcc));
defparam \delay_reg[1][1] .is_wysiwyg = "true";
defparam \delay_reg[1][1] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~30 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~30_combout ),
	.cout());
defparam \delay_reg~30 .lut_mask = 16'h8888;
defparam \delay_reg~30 .sum_lutc_input = "datac";

dffeas \delay_reg[2][1] (
	.clk(clock),
	.d(\delay_reg~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][1]~q ),
	.prn(vcc));
defparam \delay_reg[2][1] .is_wysiwyg = "true";
defparam \delay_reg[2][1] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~4 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~4_combout ),
	.cout());
defparam \delay_reg~4 .lut_mask = 16'h8888;
defparam \delay_reg~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~81 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~81_combout ),
	.cout());
defparam \delay_reg~81 .lut_mask = 16'h8888;
defparam \delay_reg~81 .sum_lutc_input = "datac";

dffeas \delay_reg[0][2] (
	.clk(clock),
	.d(\delay_reg~81_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][2]~q ),
	.prn(vcc));
defparam \delay_reg[0][2] .is_wysiwyg = "true";
defparam \delay_reg[0][2] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~57 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~57_combout ),
	.cout());
defparam \delay_reg~57 .lut_mask = 16'h8888;
defparam \delay_reg~57 .sum_lutc_input = "datac";

dffeas \delay_reg[1][2] (
	.clk(clock),
	.d(\delay_reg~57_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][2]~q ),
	.prn(vcc));
defparam \delay_reg[1][2] .is_wysiwyg = "true";
defparam \delay_reg[1][2] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~31 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~31_combout ),
	.cout());
defparam \delay_reg~31 .lut_mask = 16'h8888;
defparam \delay_reg~31 .sum_lutc_input = "datac";

dffeas \delay_reg[2][2] (
	.clk(clock),
	.d(\delay_reg~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][2]~q ),
	.prn(vcc));
defparam \delay_reg[2][2] .is_wysiwyg = "true";
defparam \delay_reg[2][2] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~5 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~5_combout ),
	.cout());
defparam \delay_reg~5 .lut_mask = 16'h8888;
defparam \delay_reg~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~82 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~82_combout ),
	.cout());
defparam \delay_reg~82 .lut_mask = 16'h8888;
defparam \delay_reg~82 .sum_lutc_input = "datac";

dffeas \delay_reg[0][3] (
	.clk(clock),
	.d(\delay_reg~82_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][3]~q ),
	.prn(vcc));
defparam \delay_reg[0][3] .is_wysiwyg = "true";
defparam \delay_reg[0][3] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~58 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~58_combout ),
	.cout());
defparam \delay_reg~58 .lut_mask = 16'h8888;
defparam \delay_reg~58 .sum_lutc_input = "datac";

dffeas \delay_reg[1][3] (
	.clk(clock),
	.d(\delay_reg~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][3]~q ),
	.prn(vcc));
defparam \delay_reg[1][3] .is_wysiwyg = "true";
defparam \delay_reg[1][3] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~32 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~32_combout ),
	.cout());
defparam \delay_reg~32 .lut_mask = 16'h8888;
defparam \delay_reg~32 .sum_lutc_input = "datac";

dffeas \delay_reg[2][3] (
	.clk(clock),
	.d(\delay_reg~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][3]~q ),
	.prn(vcc));
defparam \delay_reg[2][3] .is_wysiwyg = "true";
defparam \delay_reg[2][3] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~6 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~6_combout ),
	.cout());
defparam \delay_reg~6 .lut_mask = 16'h8888;
defparam \delay_reg~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~83 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~83_combout ),
	.cout());
defparam \delay_reg~83 .lut_mask = 16'h8888;
defparam \delay_reg~83 .sum_lutc_input = "datac";

dffeas \delay_reg[0][4] (
	.clk(clock),
	.d(\delay_reg~83_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][4]~q ),
	.prn(vcc));
defparam \delay_reg[0][4] .is_wysiwyg = "true";
defparam \delay_reg[0][4] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~59 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~59_combout ),
	.cout());
defparam \delay_reg~59 .lut_mask = 16'h8888;
defparam \delay_reg~59 .sum_lutc_input = "datac";

dffeas \delay_reg[1][4] (
	.clk(clock),
	.d(\delay_reg~59_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][4]~q ),
	.prn(vcc));
defparam \delay_reg[1][4] .is_wysiwyg = "true";
defparam \delay_reg[1][4] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~33 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~33_combout ),
	.cout());
defparam \delay_reg~33 .lut_mask = 16'h8888;
defparam \delay_reg~33 .sum_lutc_input = "datac";

dffeas \delay_reg[2][4] (
	.clk(clock),
	.d(\delay_reg~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][4]~q ),
	.prn(vcc));
defparam \delay_reg[2][4] .is_wysiwyg = "true";
defparam \delay_reg[2][4] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~7 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~7_combout ),
	.cout());
defparam \delay_reg~7 .lut_mask = 16'h8888;
defparam \delay_reg~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~84 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~84_combout ),
	.cout());
defparam \delay_reg~84 .lut_mask = 16'h8888;
defparam \delay_reg~84 .sum_lutc_input = "datac";

dffeas \delay_reg[0][5] (
	.clk(clock),
	.d(\delay_reg~84_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][5]~q ),
	.prn(vcc));
defparam \delay_reg[0][5] .is_wysiwyg = "true";
defparam \delay_reg[0][5] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~60 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~60_combout ),
	.cout());
defparam \delay_reg~60 .lut_mask = 16'h8888;
defparam \delay_reg~60 .sum_lutc_input = "datac";

dffeas \delay_reg[1][5] (
	.clk(clock),
	.d(\delay_reg~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][5]~q ),
	.prn(vcc));
defparam \delay_reg[1][5] .is_wysiwyg = "true";
defparam \delay_reg[1][5] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~34 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~34_combout ),
	.cout());
defparam \delay_reg~34 .lut_mask = 16'h8888;
defparam \delay_reg~34 .sum_lutc_input = "datac";

dffeas \delay_reg[2][5] (
	.clk(clock),
	.d(\delay_reg~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][5]~q ),
	.prn(vcc));
defparam \delay_reg[2][5] .is_wysiwyg = "true";
defparam \delay_reg[2][5] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~8 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~8_combout ),
	.cout());
defparam \delay_reg~8 .lut_mask = 16'h8888;
defparam \delay_reg~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~85 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~85_combout ),
	.cout());
defparam \delay_reg~85 .lut_mask = 16'h8888;
defparam \delay_reg~85 .sum_lutc_input = "datac";

dffeas \delay_reg[0][6] (
	.clk(clock),
	.d(\delay_reg~85_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][6]~q ),
	.prn(vcc));
defparam \delay_reg[0][6] .is_wysiwyg = "true";
defparam \delay_reg[0][6] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~61 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~61_combout ),
	.cout());
defparam \delay_reg~61 .lut_mask = 16'h8888;
defparam \delay_reg~61 .sum_lutc_input = "datac";

dffeas \delay_reg[1][6] (
	.clk(clock),
	.d(\delay_reg~61_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][6]~q ),
	.prn(vcc));
defparam \delay_reg[1][6] .is_wysiwyg = "true";
defparam \delay_reg[1][6] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~35 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~35_combout ),
	.cout());
defparam \delay_reg~35 .lut_mask = 16'h8888;
defparam \delay_reg~35 .sum_lutc_input = "datac";

dffeas \delay_reg[2][6] (
	.clk(clock),
	.d(\delay_reg~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][6]~q ),
	.prn(vcc));
defparam \delay_reg[2][6] .is_wysiwyg = "true";
defparam \delay_reg[2][6] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~9 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~9_combout ),
	.cout());
defparam \delay_reg~9 .lut_mask = 16'h8888;
defparam \delay_reg~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~86 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~86_combout ),
	.cout());
defparam \delay_reg~86 .lut_mask = 16'h8888;
defparam \delay_reg~86 .sum_lutc_input = "datac";

dffeas \delay_reg[0][7] (
	.clk(clock),
	.d(\delay_reg~86_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][7]~q ),
	.prn(vcc));
defparam \delay_reg[0][7] .is_wysiwyg = "true";
defparam \delay_reg[0][7] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~62 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~62_combout ),
	.cout());
defparam \delay_reg~62 .lut_mask = 16'h8888;
defparam \delay_reg~62 .sum_lutc_input = "datac";

dffeas \delay_reg[1][7] (
	.clk(clock),
	.d(\delay_reg~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][7]~q ),
	.prn(vcc));
defparam \delay_reg[1][7] .is_wysiwyg = "true";
defparam \delay_reg[1][7] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~36 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~36_combout ),
	.cout());
defparam \delay_reg~36 .lut_mask = 16'h8888;
defparam \delay_reg~36 .sum_lutc_input = "datac";

dffeas \delay_reg[2][7] (
	.clk(clock),
	.d(\delay_reg~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][7]~q ),
	.prn(vcc));
defparam \delay_reg[2][7] .is_wysiwyg = "true";
defparam \delay_reg[2][7] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~10 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~10_combout ),
	.cout());
defparam \delay_reg~10 .lut_mask = 16'h8888;
defparam \delay_reg~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~87 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_8),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~87_combout ),
	.cout());
defparam \delay_reg~87 .lut_mask = 16'h8888;
defparam \delay_reg~87 .sum_lutc_input = "datac";

dffeas \delay_reg[0][8] (
	.clk(clock),
	.d(\delay_reg~87_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][8]~q ),
	.prn(vcc));
defparam \delay_reg[0][8] .is_wysiwyg = "true";
defparam \delay_reg[0][8] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~63 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~63_combout ),
	.cout());
defparam \delay_reg~63 .lut_mask = 16'h8888;
defparam \delay_reg~63 .sum_lutc_input = "datac";

dffeas \delay_reg[1][8] (
	.clk(clock),
	.d(\delay_reg~63_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][8]~q ),
	.prn(vcc));
defparam \delay_reg[1][8] .is_wysiwyg = "true";
defparam \delay_reg[1][8] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~37 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~37_combout ),
	.cout());
defparam \delay_reg~37 .lut_mask = 16'h8888;
defparam \delay_reg~37 .sum_lutc_input = "datac";

dffeas \delay_reg[2][8] (
	.clk(clock),
	.d(\delay_reg~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][8]~q ),
	.prn(vcc));
defparam \delay_reg[2][8] .is_wysiwyg = "true";
defparam \delay_reg[2][8] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~11 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~11_combout ),
	.cout());
defparam \delay_reg~11 .lut_mask = 16'h8888;
defparam \delay_reg~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~88 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~88_combout ),
	.cout());
defparam \delay_reg~88 .lut_mask = 16'h8888;
defparam \delay_reg~88 .sum_lutc_input = "datac";

dffeas \delay_reg[0][9] (
	.clk(clock),
	.d(\delay_reg~88_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][9]~q ),
	.prn(vcc));
defparam \delay_reg[0][9] .is_wysiwyg = "true";
defparam \delay_reg[0][9] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~64 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~64_combout ),
	.cout());
defparam \delay_reg~64 .lut_mask = 16'h8888;
defparam \delay_reg~64 .sum_lutc_input = "datac";

dffeas \delay_reg[1][9] (
	.clk(clock),
	.d(\delay_reg~64_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][9]~q ),
	.prn(vcc));
defparam \delay_reg[1][9] .is_wysiwyg = "true";
defparam \delay_reg[1][9] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~38 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~38_combout ),
	.cout());
defparam \delay_reg~38 .lut_mask = 16'h8888;
defparam \delay_reg~38 .sum_lutc_input = "datac";

dffeas \delay_reg[2][9] (
	.clk(clock),
	.d(\delay_reg~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][9]~q ),
	.prn(vcc));
defparam \delay_reg[2][9] .is_wysiwyg = "true";
defparam \delay_reg[2][9] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~12 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~12_combout ),
	.cout());
defparam \delay_reg~12 .lut_mask = 16'h8888;
defparam \delay_reg~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~89 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_10),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~89_combout ),
	.cout());
defparam \delay_reg~89 .lut_mask = 16'h8888;
defparam \delay_reg~89 .sum_lutc_input = "datac";

dffeas \delay_reg[0][10] (
	.clk(clock),
	.d(\delay_reg~89_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][10]~q ),
	.prn(vcc));
defparam \delay_reg[0][10] .is_wysiwyg = "true";
defparam \delay_reg[0][10] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~65 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~65_combout ),
	.cout());
defparam \delay_reg~65 .lut_mask = 16'h8888;
defparam \delay_reg~65 .sum_lutc_input = "datac";

dffeas \delay_reg[1][10] (
	.clk(clock),
	.d(\delay_reg~65_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][10]~q ),
	.prn(vcc));
defparam \delay_reg[1][10] .is_wysiwyg = "true";
defparam \delay_reg[1][10] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~39 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~39_combout ),
	.cout());
defparam \delay_reg~39 .lut_mask = 16'h8888;
defparam \delay_reg~39 .sum_lutc_input = "datac";

dffeas \delay_reg[2][10] (
	.clk(clock),
	.d(\delay_reg~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][10]~q ),
	.prn(vcc));
defparam \delay_reg[2][10] .is_wysiwyg = "true";
defparam \delay_reg[2][10] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~13 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~13_combout ),
	.cout());
defparam \delay_reg~13 .lut_mask = 16'h8888;
defparam \delay_reg~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~90 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~90_combout ),
	.cout());
defparam \delay_reg~90 .lut_mask = 16'h8888;
defparam \delay_reg~90 .sum_lutc_input = "datac";

dffeas \delay_reg[0][11] (
	.clk(clock),
	.d(\delay_reg~90_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][11]~q ),
	.prn(vcc));
defparam \delay_reg[0][11] .is_wysiwyg = "true";
defparam \delay_reg[0][11] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~66 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~66_combout ),
	.cout());
defparam \delay_reg~66 .lut_mask = 16'h8888;
defparam \delay_reg~66 .sum_lutc_input = "datac";

dffeas \delay_reg[1][11] (
	.clk(clock),
	.d(\delay_reg~66_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][11]~q ),
	.prn(vcc));
defparam \delay_reg[1][11] .is_wysiwyg = "true";
defparam \delay_reg[1][11] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~40 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~40_combout ),
	.cout());
defparam \delay_reg~40 .lut_mask = 16'h8888;
defparam \delay_reg~40 .sum_lutc_input = "datac";

dffeas \delay_reg[2][11] (
	.clk(clock),
	.d(\delay_reg~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][11]~q ),
	.prn(vcc));
defparam \delay_reg[2][11] .is_wysiwyg = "true";
defparam \delay_reg[2][11] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~14 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~14_combout ),
	.cout());
defparam \delay_reg~14 .lut_mask = 16'h8888;
defparam \delay_reg~14 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~91 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_12),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~91_combout ),
	.cout());
defparam \delay_reg~91 .lut_mask = 16'h8888;
defparam \delay_reg~91 .sum_lutc_input = "datac";

dffeas \delay_reg[0][12] (
	.clk(clock),
	.d(\delay_reg~91_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][12]~q ),
	.prn(vcc));
defparam \delay_reg[0][12] .is_wysiwyg = "true";
defparam \delay_reg[0][12] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~67 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~67_combout ),
	.cout());
defparam \delay_reg~67 .lut_mask = 16'h8888;
defparam \delay_reg~67 .sum_lutc_input = "datac";

dffeas \delay_reg[1][12] (
	.clk(clock),
	.d(\delay_reg~67_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][12]~q ),
	.prn(vcc));
defparam \delay_reg[1][12] .is_wysiwyg = "true";
defparam \delay_reg[1][12] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~41 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~41_combout ),
	.cout());
defparam \delay_reg~41 .lut_mask = 16'h8888;
defparam \delay_reg~41 .sum_lutc_input = "datac";

dffeas \delay_reg[2][12] (
	.clk(clock),
	.d(\delay_reg~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][12]~q ),
	.prn(vcc));
defparam \delay_reg[2][12] .is_wysiwyg = "true";
defparam \delay_reg[2][12] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~15 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~15_combout ),
	.cout());
defparam \delay_reg~15 .lut_mask = 16'h8888;
defparam \delay_reg~15 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~92 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_13),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~92_combout ),
	.cout());
defparam \delay_reg~92 .lut_mask = 16'h8888;
defparam \delay_reg~92 .sum_lutc_input = "datac";

dffeas \delay_reg[0][13] (
	.clk(clock),
	.d(\delay_reg~92_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][13]~q ),
	.prn(vcc));
defparam \delay_reg[0][13] .is_wysiwyg = "true";
defparam \delay_reg[0][13] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~68 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~68_combout ),
	.cout());
defparam \delay_reg~68 .lut_mask = 16'h8888;
defparam \delay_reg~68 .sum_lutc_input = "datac";

dffeas \delay_reg[1][13] (
	.clk(clock),
	.d(\delay_reg~68_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][13]~q ),
	.prn(vcc));
defparam \delay_reg[1][13] .is_wysiwyg = "true";
defparam \delay_reg[1][13] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~42 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~42_combout ),
	.cout());
defparam \delay_reg~42 .lut_mask = 16'h8888;
defparam \delay_reg~42 .sum_lutc_input = "datac";

dffeas \delay_reg[2][13] (
	.clk(clock),
	.d(\delay_reg~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][13]~q ),
	.prn(vcc));
defparam \delay_reg[2][13] .is_wysiwyg = "true";
defparam \delay_reg[2][13] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~16 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~16_combout ),
	.cout());
defparam \delay_reg~16 .lut_mask = 16'h8888;
defparam \delay_reg~16 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~93 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_14),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~93_combout ),
	.cout());
defparam \delay_reg~93 .lut_mask = 16'h8888;
defparam \delay_reg~93 .sum_lutc_input = "datac";

dffeas \delay_reg[0][14] (
	.clk(clock),
	.d(\delay_reg~93_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][14]~q ),
	.prn(vcc));
defparam \delay_reg[0][14] .is_wysiwyg = "true";
defparam \delay_reg[0][14] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~69 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~69_combout ),
	.cout());
defparam \delay_reg~69 .lut_mask = 16'h8888;
defparam \delay_reg~69 .sum_lutc_input = "datac";

dffeas \delay_reg[1][14] (
	.clk(clock),
	.d(\delay_reg~69_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][14]~q ),
	.prn(vcc));
defparam \delay_reg[1][14] .is_wysiwyg = "true";
defparam \delay_reg[1][14] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~43 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~43_combout ),
	.cout());
defparam \delay_reg~43 .lut_mask = 16'h8888;
defparam \delay_reg~43 .sum_lutc_input = "datac";

dffeas \delay_reg[2][14] (
	.clk(clock),
	.d(\delay_reg~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][14]~q ),
	.prn(vcc));
defparam \delay_reg[2][14] .is_wysiwyg = "true";
defparam \delay_reg[2][14] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~17 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~17_combout ),
	.cout());
defparam \delay_reg~17 .lut_mask = 16'h8888;
defparam \delay_reg~17 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~94 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_15),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~94_combout ),
	.cout());
defparam \delay_reg~94 .lut_mask = 16'h8888;
defparam \delay_reg~94 .sum_lutc_input = "datac";

dffeas \delay_reg[0][15] (
	.clk(clock),
	.d(\delay_reg~94_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][15]~q ),
	.prn(vcc));
defparam \delay_reg[0][15] .is_wysiwyg = "true";
defparam \delay_reg[0][15] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~70 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~70_combout ),
	.cout());
defparam \delay_reg~70 .lut_mask = 16'h8888;
defparam \delay_reg~70 .sum_lutc_input = "datac";

dffeas \delay_reg[1][15] (
	.clk(clock),
	.d(\delay_reg~70_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][15]~q ),
	.prn(vcc));
defparam \delay_reg[1][15] .is_wysiwyg = "true";
defparam \delay_reg[1][15] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~44 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~44_combout ),
	.cout());
defparam \delay_reg~44 .lut_mask = 16'h8888;
defparam \delay_reg~44 .sum_lutc_input = "datac";

dffeas \delay_reg[2][15] (
	.clk(clock),
	.d(\delay_reg~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][15]~q ),
	.prn(vcc));
defparam \delay_reg[2][15] .is_wysiwyg = "true";
defparam \delay_reg[2][15] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~18 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~18_combout ),
	.cout());
defparam \delay_reg~18 .lut_mask = 16'h8888;
defparam \delay_reg~18 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~95 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_16),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~95_combout ),
	.cout());
defparam \delay_reg~95 .lut_mask = 16'h8888;
defparam \delay_reg~95 .sum_lutc_input = "datac";

dffeas \delay_reg[0][16] (
	.clk(clock),
	.d(\delay_reg~95_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][16]~q ),
	.prn(vcc));
defparam \delay_reg[0][16] .is_wysiwyg = "true";
defparam \delay_reg[0][16] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~71 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~71_combout ),
	.cout());
defparam \delay_reg~71 .lut_mask = 16'h8888;
defparam \delay_reg~71 .sum_lutc_input = "datac";

dffeas \delay_reg[1][16] (
	.clk(clock),
	.d(\delay_reg~71_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][16]~q ),
	.prn(vcc));
defparam \delay_reg[1][16] .is_wysiwyg = "true";
defparam \delay_reg[1][16] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~45 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~45_combout ),
	.cout());
defparam \delay_reg~45 .lut_mask = 16'h8888;
defparam \delay_reg~45 .sum_lutc_input = "datac";

dffeas \delay_reg[2][16] (
	.clk(clock),
	.d(\delay_reg~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][16]~q ),
	.prn(vcc));
defparam \delay_reg[2][16] .is_wysiwyg = "true";
defparam \delay_reg[2][16] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~19 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~19_combout ),
	.cout());
defparam \delay_reg~19 .lut_mask = 16'h8888;
defparam \delay_reg~19 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~96 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_17),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~96_combout ),
	.cout());
defparam \delay_reg~96 .lut_mask = 16'h8888;
defparam \delay_reg~96 .sum_lutc_input = "datac";

dffeas \delay_reg[0][17] (
	.clk(clock),
	.d(\delay_reg~96_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][17]~q ),
	.prn(vcc));
defparam \delay_reg[0][17] .is_wysiwyg = "true";
defparam \delay_reg[0][17] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~72 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][17]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~72_combout ),
	.cout());
defparam \delay_reg~72 .lut_mask = 16'h8888;
defparam \delay_reg~72 .sum_lutc_input = "datac";

dffeas \delay_reg[1][17] (
	.clk(clock),
	.d(\delay_reg~72_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][17]~q ),
	.prn(vcc));
defparam \delay_reg[1][17] .is_wysiwyg = "true";
defparam \delay_reg[1][17] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~46 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][17]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~46_combout ),
	.cout());
defparam \delay_reg~46 .lut_mask = 16'h8888;
defparam \delay_reg~46 .sum_lutc_input = "datac";

dffeas \delay_reg[2][17] (
	.clk(clock),
	.d(\delay_reg~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][17]~q ),
	.prn(vcc));
defparam \delay_reg[2][17] .is_wysiwyg = "true";
defparam \delay_reg[2][17] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~20 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][17]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~20_combout ),
	.cout());
defparam \delay_reg~20 .lut_mask = 16'h8888;
defparam \delay_reg~20 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~97 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_18),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~97_combout ),
	.cout());
defparam \delay_reg~97 .lut_mask = 16'h8888;
defparam \delay_reg~97 .sum_lutc_input = "datac";

dffeas \delay_reg[0][18] (
	.clk(clock),
	.d(\delay_reg~97_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][18]~q ),
	.prn(vcc));
defparam \delay_reg[0][18] .is_wysiwyg = "true";
defparam \delay_reg[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~73 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][18]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~73_combout ),
	.cout());
defparam \delay_reg~73 .lut_mask = 16'h8888;
defparam \delay_reg~73 .sum_lutc_input = "datac";

dffeas \delay_reg[1][18] (
	.clk(clock),
	.d(\delay_reg~73_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][18]~q ),
	.prn(vcc));
defparam \delay_reg[1][18] .is_wysiwyg = "true";
defparam \delay_reg[1][18] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~47 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][18]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~47_combout ),
	.cout());
defparam \delay_reg~47 .lut_mask = 16'h8888;
defparam \delay_reg~47 .sum_lutc_input = "datac";

dffeas \delay_reg[2][18] (
	.clk(clock),
	.d(\delay_reg~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][18]~q ),
	.prn(vcc));
defparam \delay_reg[2][18] .is_wysiwyg = "true";
defparam \delay_reg[2][18] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~21 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][18]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~21_combout ),
	.cout());
defparam \delay_reg~21 .lut_mask = 16'h8888;
defparam \delay_reg~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~98 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_19),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~98_combout ),
	.cout());
defparam \delay_reg~98 .lut_mask = 16'h8888;
defparam \delay_reg~98 .sum_lutc_input = "datac";

dffeas \delay_reg[0][19] (
	.clk(clock),
	.d(\delay_reg~98_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][19]~q ),
	.prn(vcc));
defparam \delay_reg[0][19] .is_wysiwyg = "true";
defparam \delay_reg[0][19] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~74 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][19]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~74_combout ),
	.cout());
defparam \delay_reg~74 .lut_mask = 16'h8888;
defparam \delay_reg~74 .sum_lutc_input = "datac";

dffeas \delay_reg[1][19] (
	.clk(clock),
	.d(\delay_reg~74_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][19]~q ),
	.prn(vcc));
defparam \delay_reg[1][19] .is_wysiwyg = "true";
defparam \delay_reg[1][19] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~48 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][19]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~48_combout ),
	.cout());
defparam \delay_reg~48 .lut_mask = 16'h8888;
defparam \delay_reg~48 .sum_lutc_input = "datac";

dffeas \delay_reg[2][19] (
	.clk(clock),
	.d(\delay_reg~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][19]~q ),
	.prn(vcc));
defparam \delay_reg[2][19] .is_wysiwyg = "true";
defparam \delay_reg[2][19] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~22 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][19]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~22_combout ),
	.cout());
defparam \delay_reg~22 .lut_mask = 16'h8888;
defparam \delay_reg~22 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~99 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_20),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~99_combout ),
	.cout());
defparam \delay_reg~99 .lut_mask = 16'h8888;
defparam \delay_reg~99 .sum_lutc_input = "datac";

dffeas \delay_reg[0][20] (
	.clk(clock),
	.d(\delay_reg~99_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][20]~q ),
	.prn(vcc));
defparam \delay_reg[0][20] .is_wysiwyg = "true";
defparam \delay_reg[0][20] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~75 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~75_combout ),
	.cout());
defparam \delay_reg~75 .lut_mask = 16'h8888;
defparam \delay_reg~75 .sum_lutc_input = "datac";

dffeas \delay_reg[1][20] (
	.clk(clock),
	.d(\delay_reg~75_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][20]~q ),
	.prn(vcc));
defparam \delay_reg[1][20] .is_wysiwyg = "true";
defparam \delay_reg[1][20] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~49 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~49_combout ),
	.cout());
defparam \delay_reg~49 .lut_mask = 16'h8888;
defparam \delay_reg~49 .sum_lutc_input = "datac";

dffeas \delay_reg[2][20] (
	.clk(clock),
	.d(\delay_reg~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][20]~q ),
	.prn(vcc));
defparam \delay_reg[2][20] .is_wysiwyg = "true";
defparam \delay_reg[2][20] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~23 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~23_combout ),
	.cout());
defparam \delay_reg~23 .lut_mask = 16'h8888;
defparam \delay_reg~23 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~100 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_21),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~100_combout ),
	.cout());
defparam \delay_reg~100 .lut_mask = 16'h8888;
defparam \delay_reg~100 .sum_lutc_input = "datac";

dffeas \delay_reg[0][21] (
	.clk(clock),
	.d(\delay_reg~100_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][21]~q ),
	.prn(vcc));
defparam \delay_reg[0][21] .is_wysiwyg = "true";
defparam \delay_reg[0][21] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~76 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][21]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~76_combout ),
	.cout());
defparam \delay_reg~76 .lut_mask = 16'h8888;
defparam \delay_reg~76 .sum_lutc_input = "datac";

dffeas \delay_reg[1][21] (
	.clk(clock),
	.d(\delay_reg~76_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][21]~q ),
	.prn(vcc));
defparam \delay_reg[1][21] .is_wysiwyg = "true";
defparam \delay_reg[1][21] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~50 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][21]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~50_combout ),
	.cout());
defparam \delay_reg~50 .lut_mask = 16'h8888;
defparam \delay_reg~50 .sum_lutc_input = "datac";

dffeas \delay_reg[2][21] (
	.clk(clock),
	.d(\delay_reg~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][21]~q ),
	.prn(vcc));
defparam \delay_reg[2][21] .is_wysiwyg = "true";
defparam \delay_reg[2][21] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~24 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][21]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~24_combout ),
	.cout());
defparam \delay_reg~24 .lut_mask = 16'h8888;
defparam \delay_reg~24 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~101 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_22),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~101_combout ),
	.cout());
defparam \delay_reg~101 .lut_mask = 16'h8888;
defparam \delay_reg~101 .sum_lutc_input = "datac";

dffeas \delay_reg[0][22] (
	.clk(clock),
	.d(\delay_reg~101_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][22]~q ),
	.prn(vcc));
defparam \delay_reg[0][22] .is_wysiwyg = "true";
defparam \delay_reg[0][22] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~77 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][22]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~77_combout ),
	.cout());
defparam \delay_reg~77 .lut_mask = 16'h8888;
defparam \delay_reg~77 .sum_lutc_input = "datac";

dffeas \delay_reg[1][22] (
	.clk(clock),
	.d(\delay_reg~77_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][22]~q ),
	.prn(vcc));
defparam \delay_reg[1][22] .is_wysiwyg = "true";
defparam \delay_reg[1][22] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~51 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][22]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~51_combout ),
	.cout());
defparam \delay_reg~51 .lut_mask = 16'h8888;
defparam \delay_reg~51 .sum_lutc_input = "datac";

dffeas \delay_reg[2][22] (
	.clk(clock),
	.d(\delay_reg~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][22]~q ),
	.prn(vcc));
defparam \delay_reg[2][22] .is_wysiwyg = "true";
defparam \delay_reg[2][22] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~25 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][22]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~25_combout ),
	.cout());
defparam \delay_reg~25 .lut_mask = 16'h8888;
defparam \delay_reg~25 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~102 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(data_out_23),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~102_combout ),
	.cout());
defparam \delay_reg~102 .lut_mask = 16'h8888;
defparam \delay_reg~102 .sum_lutc_input = "datac";

dffeas \delay_reg[0][23] (
	.clk(clock),
	.d(\delay_reg~102_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[0][23]~q ),
	.prn(vcc));
defparam \delay_reg[0][23] .is_wysiwyg = "true";
defparam \delay_reg[0][23] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~78 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[0][23]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~78_combout ),
	.cout());
defparam \delay_reg~78 .lut_mask = 16'h8888;
defparam \delay_reg~78 .sum_lutc_input = "datac";

dffeas \delay_reg[1][23] (
	.clk(clock),
	.d(\delay_reg~78_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[1][23]~q ),
	.prn(vcc));
defparam \delay_reg[1][23] .is_wysiwyg = "true";
defparam \delay_reg[1][23] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~52 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[1][23]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~52_combout ),
	.cout());
defparam \delay_reg~52 .lut_mask = 16'h8888;
defparam \delay_reg~52 .sum_lutc_input = "datac";

dffeas \delay_reg[2][23] (
	.clk(clock),
	.d(\delay_reg~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][23]~q ),
	.prn(vcc));
defparam \delay_reg[2][23] .is_wysiwyg = "true";
defparam \delay_reg[2][23] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~26 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][23]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~26_combout ),
	.cout());
defparam \delay_reg~26 .lut_mask = 16'h8888;
defparam \delay_reg~26 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \delay_reg~53 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(delay_reg_24_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~53_combout ),
	.cout());
defparam \delay_reg~53 .lut_mask = 16'h8888;
defparam \delay_reg~53 .sum_lutc_input = "datac";

dffeas \delay_reg[2][24] (
	.clk(clock),
	.d(\delay_reg~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delay_reg[2][24]~q ),
	.prn(vcc));
defparam \delay_reg[2][24] .is_wysiwyg = "true";
defparam \delay_reg[2][24] .power_up = "low";

fiftyfivenm_lcell_comb \delay_reg~27 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\delay_reg[2][24]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_reg~27_combout ),
	.cout());
defparam \delay_reg~27 .lut_mask = 16'h8888;
defparam \delay_reg~27 .sum_lutc_input = "datac";

endmodule

module lms_dsp_dual_running_sum (
	short_sum_reg_0,
	short_sum_reg_1,
	short_sum_reg_2,
	short_sum_reg_3,
	short_sum_reg_4,
	short_sum_reg_5,
	short_sum_reg_6,
	short_sum_reg_7,
	short_sum_reg_8,
	short_sum_reg_9,
	short_sum_reg_10,
	short_sum_reg_11,
	short_sum_reg_12,
	short_sum_reg_13,
	short_sum_reg_14,
	short_sum_reg_15,
	short_sum_reg_16,
	short_sum_reg_17,
	LessThan0,
	mag_reg_0,
	running_reg,
	mag_reg_1,
	mag_reg_2,
	mag_reg_3,
	mag_reg_4,
	mag_reg_5,
	mag_reg_6,
	mag_reg_7,
	mag_reg_8,
	mag_reg_9,
	mag_reg_10,
	mag_reg_11,
	mag_reg_12,
	long_shift_rescale_0,
	long_shift_rescale_1,
	long_shift_rescale_2,
	long_shift_rescale_3,
	long_shift_rescale_4,
	long_shift_rescale_5,
	long_shift_rescale_6,
	long_shift_rescale_7,
	long_shift_rescale_8,
	long_shift_rescale_9,
	long_shift_rescale_10,
	long_shift_rescale_11,
	long_shift_rescale_12,
	long_shift_rescale_13,
	long_shift_rescale_14,
	long_shift_rescale_15,
	long_shift_rescale_16,
	long_shift_rescale_17,
	long_shift_rescale_18,
	long_shift_rescale_19,
	long_shift_rescale_20,
	altera_reset_synchronizer_int_chain_out,
	launch1,
	long_shift_rescale_25,
	launch2,
	delay_reg_24_0,
	GND_port,
	clk_clk,
	ppd_cfg_clear_rs,
	ppd_cfg_threshold_0,
	ppd_cfg_threshold_1,
	ppd_cfg_threshold_2,
	ppd_cfg_threshold_3,
	ppd_cfg_threshold_4,
	ppd_cfg_threshold_5,
	ppd_cfg_threshold_6,
	ppd_cfg_threshold_7)/* synthesis synthesis_greybox=0 */;
output 	short_sum_reg_0;
output 	short_sum_reg_1;
output 	short_sum_reg_2;
output 	short_sum_reg_3;
output 	short_sum_reg_4;
output 	short_sum_reg_5;
output 	short_sum_reg_6;
output 	short_sum_reg_7;
output 	short_sum_reg_8;
output 	short_sum_reg_9;
output 	short_sum_reg_10;
output 	short_sum_reg_11;
output 	short_sum_reg_12;
output 	short_sum_reg_13;
output 	short_sum_reg_14;
output 	short_sum_reg_15;
output 	short_sum_reg_16;
output 	short_sum_reg_17;
output 	LessThan0;
input 	mag_reg_0;
input 	running_reg;
input 	mag_reg_1;
input 	mag_reg_2;
input 	mag_reg_3;
input 	mag_reg_4;
input 	mag_reg_5;
input 	mag_reg_6;
input 	mag_reg_7;
input 	mag_reg_8;
input 	mag_reg_9;
input 	mag_reg_10;
input 	mag_reg_11;
input 	mag_reg_12;
output 	long_shift_rescale_0;
output 	long_shift_rescale_1;
output 	long_shift_rescale_2;
output 	long_shift_rescale_3;
output 	long_shift_rescale_4;
output 	long_shift_rescale_5;
output 	long_shift_rescale_6;
output 	long_shift_rescale_7;
output 	long_shift_rescale_8;
output 	long_shift_rescale_9;
output 	long_shift_rescale_10;
output 	long_shift_rescale_11;
output 	long_shift_rescale_12;
output 	long_shift_rescale_13;
output 	long_shift_rescale_14;
output 	long_shift_rescale_15;
output 	long_shift_rescale_16;
output 	long_shift_rescale_17;
output 	long_shift_rescale_18;
output 	long_shift_rescale_19;
output 	long_shift_rescale_20;
input 	altera_reset_synchronizer_int_chain_out;
output 	launch1;
output 	long_shift_rescale_25;
output 	launch2;
input 	delay_reg_24_0;
input 	GND_port;
input 	clk_clk;
input 	ppd_cfg_clear_rs;
input 	ppd_cfg_threshold_0;
input 	ppd_cfg_threshold_1;
input 	ppd_cfg_threshold_2;
input 	ppd_cfg_threshold_3;
input 	ppd_cfg_threshold_4;
input 	ppd_cfg_threshold_5;
input 	ppd_cfg_threshold_6;
input 	ppd_cfg_threshold_7;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mult0|auto_generated|w138w[0] ;
wire \Mult0|auto_generated|w138w[1] ;
wire \Mult0|auto_generated|w138w[2] ;
wire \short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[0] ;
wire \short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[1] ;
wire \short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[2] ;
wire \short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[3] ;
wire \short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[4] ;
wire \short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[5] ;
wire \short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[6] ;
wire \short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[7] ;
wire \short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[8] ;
wire \short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[9] ;
wire \short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[10] ;
wire \short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[11] ;
wire \short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[12] ;
wire \short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[13] ;
wire \short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[14] ;
wire \short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[15] ;
wire \long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[0] ;
wire \long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[1] ;
wire \long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[2] ;
wire \long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[3] ;
wire \long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[4] ;
wire \long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[5] ;
wire \long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[6] ;
wire \long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[7] ;
wire \long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[8] ;
wire \long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[9] ;
wire \long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[10] ;
wire \long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[11] ;
wire \long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[12] ;
wire \long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[13] ;
wire \long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[14] ;
wire \long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[15] ;
wire \Add0~0_combout ;
wire \short_sum_reg[0]~18_combout ;
wire \always0~1_combout ;
wire \always0~2_combout ;
wire \short_sum_reg[11]~20_combout ;
wire \Add0~1 ;
wire \Add0~2_combout ;
wire \short_sum_reg[0]~19 ;
wire \short_sum_reg[1]~21_combout ;
wire \Add0~3 ;
wire \Add0~4_combout ;
wire \short_sum_reg[1]~22 ;
wire \short_sum_reg[2]~23_combout ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \short_sum_reg[2]~24 ;
wire \short_sum_reg[3]~25_combout ;
wire \Add0~7 ;
wire \Add0~8_combout ;
wire \short_sum_reg[3]~26 ;
wire \short_sum_reg[4]~27_combout ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \short_sum_reg[4]~28 ;
wire \short_sum_reg[5]~29_combout ;
wire \Add0~11 ;
wire \Add0~12_combout ;
wire \short_sum_reg[5]~30 ;
wire \short_sum_reg[6]~31_combout ;
wire \Add0~13 ;
wire \Add0~14_combout ;
wire \short_sum_reg[6]~32 ;
wire \short_sum_reg[7]~33_combout ;
wire \Add0~15 ;
wire \Add0~16_combout ;
wire \short_sum_reg[7]~34 ;
wire \short_sum_reg[8]~35_combout ;
wire \Add0~17 ;
wire \Add0~18_combout ;
wire \short_sum_reg[8]~36 ;
wire \short_sum_reg[9]~37_combout ;
wire \Add0~19 ;
wire \Add0~20_combout ;
wire \short_sum_reg[9]~38 ;
wire \short_sum_reg[10]~39_combout ;
wire \Add0~21 ;
wire \Add0~22_combout ;
wire \short_sum_reg[10]~40 ;
wire \short_sum_reg[11]~41_combout ;
wire \Add0~23 ;
wire \Add0~24_combout ;
wire \short_sum_reg[11]~42 ;
wire \short_sum_reg[12]~43_combout ;
wire \Add0~25 ;
wire \Add0~26_combout ;
wire \short_sum_reg[12]~44 ;
wire \short_sum_reg[13]~45_combout ;
wire \Add0~27 ;
wire \Add0~28_combout ;
wire \short_sum_reg[13]~46 ;
wire \short_sum_reg[14]~47_combout ;
wire \Add0~29 ;
wire \Add0~30_combout ;
wire \short_sum_reg[14]~48 ;
wire \short_sum_reg[15]~49_combout ;
wire \Add0~31 ;
wire \Add0~32_combout ;
wire \short_sum_reg[15]~50 ;
wire \short_sum_reg[16]~51_combout ;
wire \Add0~33 ;
wire \Add0~34_combout ;
wire \short_sum_reg[16]~52 ;
wire \short_sum_reg[17]~53_combout ;
wire \LessThan0~1_cout ;
wire \LessThan0~3_cout ;
wire \LessThan0~5_cout ;
wire \LessThan0~7_cout ;
wire \LessThan0~9_cout ;
wire \LessThan0~11_cout ;
wire \LessThan0~13_cout ;
wire \LessThan0~15_cout ;
wire \LessThan0~17_cout ;
wire \LessThan0~19_cout ;
wire \LessThan0~21_cout ;
wire \LessThan0~23_cout ;
wire \LessThan0~25_cout ;
wire \LessThan0~27_cout ;
wire \LessThan0~29_cout ;
wire \LessThan0~31_cout ;
wire \LessThan0~33_cout ;
wire \Add3~0_combout ;
wire \long_sum_reg[0]~21_combout ;
wire \always0~0_combout ;
wire \short_counter[0]~5_combout ;
wire \short_to_long_arrived~0_combout ;
wire \short_to_long_arrived~1_combout ;
wire \short_to_long_arrived~q ;
wire \short_counter[0]~15_combout ;
wire \short_counter[0]~16_combout ;
wire \short_counter[0]~17_combout ;
wire \short_counter[0]~q ;
wire \short_counter[0]~6 ;
wire \short_counter[1]~7_combout ;
wire \short_counter[1]~q ;
wire \short_counter[1]~8 ;
wire \short_counter[2]~9_combout ;
wire \short_counter[2]~q ;
wire \short_counter[2]~10 ;
wire \short_counter[3]~11_combout ;
wire \short_counter[3]~q ;
wire \short_counter[3]~12 ;
wire \short_counter[4]~13_combout ;
wire \short_counter[4]~q ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \short_shift_full~0_combout ;
wire \short_shift_full~q ;
wire \long_sum_reg[1]~23_combout ;
wire \long_sum_reg[0]~q ;
wire \Add3~1 ;
wire \Add3~2_combout ;
wire \long_sum_reg[0]~22 ;
wire \long_sum_reg[1]~24_combout ;
wire \long_sum_reg[1]~q ;
wire \Add3~3 ;
wire \Add3~4_combout ;
wire \long_sum_reg[1]~25 ;
wire \long_sum_reg[2]~26_combout ;
wire \long_sum_reg[2]~q ;
wire \Add3~5 ;
wire \Add3~6_combout ;
wire \long_sum_reg[2]~27 ;
wire \long_sum_reg[3]~28_combout ;
wire \long_sum_reg[3]~q ;
wire \Add3~7 ;
wire \Add3~8_combout ;
wire \long_sum_reg[3]~29 ;
wire \long_sum_reg[4]~30_combout ;
wire \long_sum_reg[4]~q ;
wire \Add3~9 ;
wire \Add3~10_combout ;
wire \long_sum_reg[4]~31 ;
wire \long_sum_reg[5]~32_combout ;
wire \long_sum_reg[5]~q ;
wire \Add3~11 ;
wire \Add3~12_combout ;
wire \long_sum_reg[5]~33 ;
wire \long_sum_reg[6]~34_combout ;
wire \long_sum_reg[6]~q ;
wire \Add3~13 ;
wire \Add3~14_combout ;
wire \long_sum_reg[6]~35 ;
wire \long_sum_reg[7]~36_combout ;
wire \long_sum_reg[7]~q ;
wire \Add3~15 ;
wire \Add3~16_combout ;
wire \long_sum_reg[7]~37 ;
wire \long_sum_reg[8]~38_combout ;
wire \long_sum_reg[8]~q ;
wire \Add3~17 ;
wire \Add3~18_combout ;
wire \long_sum_reg[8]~39 ;
wire \long_sum_reg[9]~40_combout ;
wire \long_sum_reg[9]~q ;
wire \Add3~19 ;
wire \Add3~20_combout ;
wire \long_sum_reg[9]~41 ;
wire \long_sum_reg[10]~42_combout ;
wire \long_sum_reg[10]~q ;
wire \Add3~21 ;
wire \Add3~22_combout ;
wire \long_sum_reg[10]~43 ;
wire \long_sum_reg[11]~44_combout ;
wire \long_sum_reg[11]~q ;
wire \Add3~23 ;
wire \Add3~24_combout ;
wire \long_sum_reg[11]~45 ;
wire \long_sum_reg[12]~46_combout ;
wire \long_sum_reg[12]~q ;
wire \Add3~25 ;
wire \Add3~26_combout ;
wire \long_sum_reg[12]~47 ;
wire \long_sum_reg[13]~48_combout ;
wire \long_sum_reg[13]~q ;
wire \Add3~27 ;
wire \Add3~28_combout ;
wire \long_sum_reg[13]~49 ;
wire \long_sum_reg[14]~50_combout ;
wire \long_sum_reg[14]~q ;
wire \Add3~29 ;
wire \Add3~30_combout ;
wire \long_sum_reg[14]~51 ;
wire \long_sum_reg[15]~52_combout ;
wire \long_sum_reg[15]~q ;
wire \Add3~31 ;
wire \Add3~32_combout ;
wire \long_sum_reg[15]~53 ;
wire \long_sum_reg[16]~54_combout ;
wire \long_sum_reg[16]~q ;
wire \Add3~33 ;
wire \Add3~34_combout ;
wire \long_sum_reg[16]~55 ;
wire \long_sum_reg[17]~56_combout ;
wire \long_sum_reg[17]~q ;
wire \Mult0|auto_generated|mac_mult1~dataout ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT1 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT2 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT3 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT4 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT5 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT6 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT7 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT8 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT9 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT10 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT11 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT12 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT13 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT14 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT15 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT16 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT17 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT18 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT19 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT20 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT21 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT22 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT23 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT24 ;
wire \Mult0|auto_generated|mac_mult1~DATAOUT25 ;
wire \Mult0|auto_generated|w138w[3] ;
wire \long_shift_rescale~22_combout ;
wire \Mult0|auto_generated|w138w[4] ;
wire \long_shift_rescale~23_combout ;
wire \Mult0|auto_generated|w138w[5] ;
wire \long_shift_rescale~24_combout ;
wire \Mult0|auto_generated|w138w[6] ;
wire \long_shift_rescale~25_combout ;
wire \Mult0|auto_generated|w138w[7] ;
wire \long_shift_rescale~26_combout ;
wire \Mult0|auto_generated|w138w[8] ;
wire \long_shift_rescale~27_combout ;
wire \Mult0|auto_generated|w138w[9] ;
wire \long_shift_rescale~28_combout ;
wire \Mult0|auto_generated|w138w[10] ;
wire \long_shift_rescale~29_combout ;
wire \Mult0|auto_generated|w138w[11] ;
wire \long_shift_rescale~30_combout ;
wire \Mult0|auto_generated|w138w[12] ;
wire \long_shift_rescale~31_combout ;
wire \Mult0|auto_generated|w138w[13] ;
wire \long_shift_rescale~32_combout ;
wire \Mult0|auto_generated|w138w[14] ;
wire \long_shift_rescale~33_combout ;
wire \Mult0|auto_generated|w138w[15] ;
wire \long_shift_rescale~34_combout ;
wire \Mult0|auto_generated|w138w[16] ;
wire \long_shift_rescale~35_combout ;
wire \Mult0|auto_generated|w138w[17] ;
wire \long_shift_rescale~36_combout ;
wire \Add3~35 ;
wire \Add3~36_combout ;
wire \long_sum_reg[17]~57 ;
wire \long_sum_reg[18]~58_combout ;
wire \long_sum_reg[18]~q ;
wire \Add3~37 ;
wire \Add3~38_combout ;
wire \long_sum_reg[18]~59 ;
wire \long_sum_reg[19]~60_combout ;
wire \long_sum_reg[19]~q ;
wire \Add3~39 ;
wire \Add3~40_combout ;
wire \long_sum_reg[19]~61 ;
wire \long_sum_reg[20]~62_combout ;
wire \long_sum_reg[20]~q ;
wire \Mult0|auto_generated|mac_mult3~dataout ;
wire \Mult0|auto_generated|mac_mult3~DATAOUT1 ;
wire \Mult0|auto_generated|mac_mult3~DATAOUT2 ;
wire \Mult0|auto_generated|mac_mult3~DATAOUT3 ;
wire \Mult0|auto_generated|mac_mult3~DATAOUT4 ;
wire \Mult0|auto_generated|mac_mult3~DATAOUT5 ;
wire \Mult0|auto_generated|mac_mult3~DATAOUT6 ;
wire \Mult0|auto_generated|mac_mult3~DATAOUT7 ;
wire \Mult0|auto_generated|mac_mult3~DATAOUT8 ;
wire \Mult0|auto_generated|mac_mult3~DATAOUT9 ;
wire \Mult0|auto_generated|mac_mult3~DATAOUT10 ;
wire \Mult0|auto_generated|mac_out4~dataout ;
wire \Mult0|auto_generated|mac_out2~DATAOUT18 ;
wire \Mult0|auto_generated|op_1~0_combout ;
wire \long_shift_rescale~37_combout ;
wire \Mult0|auto_generated|mac_out4~DATAOUT1 ;
wire \Mult0|auto_generated|mac_out2~DATAOUT19 ;
wire \Mult0|auto_generated|op_1~1 ;
wire \Mult0|auto_generated|op_1~2_combout ;
wire \long_shift_rescale~38_combout ;
wire \Mult0|auto_generated|mac_out4~DATAOUT2 ;
wire \Mult0|auto_generated|mac_out2~DATAOUT20 ;
wire \Mult0|auto_generated|op_1~3 ;
wire \Mult0|auto_generated|op_1~4_combout ;
wire \long_shift_rescale~39_combout ;
wire \Mult0|auto_generated|mac_out4~DATAOUT3 ;
wire \Mult0|auto_generated|mac_out2~DATAOUT21 ;
wire \Mult0|auto_generated|op_1~5 ;
wire \Mult0|auto_generated|op_1~6_combout ;
wire \long_shift_rescale~40_combout ;
wire \Mult0|auto_generated|mac_out4~DATAOUT4 ;
wire \Mult0|auto_generated|mac_out2~DATAOUT22 ;
wire \Mult0|auto_generated|op_1~7 ;
wire \Mult0|auto_generated|op_1~8_combout ;
wire \long_shift_rescale~41_combout ;
wire \Mult0|auto_generated|mac_out4~DATAOUT5 ;
wire \Mult0|auto_generated|mac_out2~DATAOUT23 ;
wire \Mult0|auto_generated|op_1~9 ;
wire \Mult0|auto_generated|op_1~10_combout ;
wire \long_shift_rescale~42_combout ;
wire \long_counter[0]~8_combout ;
wire \long_counter[0]~9 ;
wire \long_counter[1]~11_combout ;
wire \long_counter[1]~q ;
wire \long_counter[1]~12 ;
wire \long_counter[2]~13_combout ;
wire \long_counter[2]~q ;
wire \long_counter[2]~14 ;
wire \long_counter[3]~15_combout ;
wire \long_counter[3]~q ;
wire \long_counter[3]~16 ;
wire \long_counter[4]~17_combout ;
wire \long_counter[4]~q ;
wire \long_counter[4]~18 ;
wire \long_counter[5]~19_combout ;
wire \long_counter[5]~q ;
wire \long_counter[5]~20 ;
wire \long_counter[6]~21_combout ;
wire \long_counter[6]~q ;
wire \long_counter[6]~22 ;
wire \long_counter[7]~23_combout ;
wire \long_counter[7]~q ;
wire \Equal1~1_combout ;
wire \long_counter[0]~10_combout ;
wire \long_counter[0]~q ;
wire \Equal1~0_combout ;
wire \launch~0_combout ;
wire \Mult0|auto_generated|mac_out4~DATAOUT6 ;
wire \Mult0|auto_generated|mac_out2~DATAOUT24 ;
wire \Mult0|auto_generated|op_1~11 ;
wire \Mult0|auto_generated|op_1~12_combout ;
wire \long_shift_rescale~43_combout ;
wire \long_shift_rescale[21]~q ;
wire \Mult0|auto_generated|mac_out4~DATAOUT7 ;
wire \Mult0|auto_generated|mac_out2~DATAOUT25 ;
wire \Mult0|auto_generated|op_1~13 ;
wire \Mult0|auto_generated|op_1~14_combout ;
wire \long_shift_rescale~44_combout ;
wire \long_shift_rescale[22]~q ;
wire \Mult0|auto_generated|mac_out4~DATAOUT8 ;
wire \Mult0|auto_generated|op_1~15 ;
wire \Mult0|auto_generated|op_1~16_combout ;
wire \long_shift_rescale~45_combout ;
wire \long_shift_rescale[23]~q ;
wire \Mult0|auto_generated|mac_out4~DATAOUT9 ;
wire \Mult0|auto_generated|op_1~17 ;
wire \Mult0|auto_generated|op_1~18_combout ;
wire \long_shift_rescale~46_combout ;
wire \long_shift_rescale[24]~q ;
wire \launch~1_combout ;
wire \Mult0|auto_generated|mac_out4~DATAOUT10 ;
wire \Mult0|auto_generated|op_1~19 ;
wire \Mult0|auto_generated|op_1~20_combout ;
wire \long_shift_rescale~47_combout ;

wire [35:0] \Mult0|auto_generated|mac_out2_DATAOUT_bus ;
wire [35:0] \Mult0|auto_generated|mac_out4_DATAOUT_bus ;
wire [35:0] \Mult0|auto_generated|mac_mult1_DATAOUT_bus ;
wire [35:0] \Mult0|auto_generated|mac_mult3_DATAOUT_bus ;

assign \Mult0|auto_generated|w138w[0]  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [0];
assign \Mult0|auto_generated|w138w[1]  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [1];
assign \Mult0|auto_generated|w138w[2]  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [2];
assign \Mult0|auto_generated|w138w[3]  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [3];
assign \Mult0|auto_generated|w138w[4]  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [4];
assign \Mult0|auto_generated|w138w[5]  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [5];
assign \Mult0|auto_generated|w138w[6]  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [6];
assign \Mult0|auto_generated|w138w[7]  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [7];
assign \Mult0|auto_generated|w138w[8]  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [8];
assign \Mult0|auto_generated|w138w[9]  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [9];
assign \Mult0|auto_generated|w138w[10]  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [10];
assign \Mult0|auto_generated|w138w[11]  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [11];
assign \Mult0|auto_generated|w138w[12]  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [12];
assign \Mult0|auto_generated|w138w[13]  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [13];
assign \Mult0|auto_generated|w138w[14]  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [14];
assign \Mult0|auto_generated|w138w[15]  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [15];
assign \Mult0|auto_generated|w138w[16]  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [16];
assign \Mult0|auto_generated|w138w[17]  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [17];
assign \Mult0|auto_generated|mac_out2~DATAOUT18  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [18];
assign \Mult0|auto_generated|mac_out2~DATAOUT19  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [19];
assign \Mult0|auto_generated|mac_out2~DATAOUT20  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [20];
assign \Mult0|auto_generated|mac_out2~DATAOUT21  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [21];
assign \Mult0|auto_generated|mac_out2~DATAOUT22  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [22];
assign \Mult0|auto_generated|mac_out2~DATAOUT23  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [23];
assign \Mult0|auto_generated|mac_out2~DATAOUT24  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [24];
assign \Mult0|auto_generated|mac_out2~DATAOUT25  = \Mult0|auto_generated|mac_out2_DATAOUT_bus [25];

assign \Mult0|auto_generated|mac_out4~dataout  = \Mult0|auto_generated|mac_out4_DATAOUT_bus [0];
assign \Mult0|auto_generated|mac_out4~DATAOUT1  = \Mult0|auto_generated|mac_out4_DATAOUT_bus [1];
assign \Mult0|auto_generated|mac_out4~DATAOUT2  = \Mult0|auto_generated|mac_out4_DATAOUT_bus [2];
assign \Mult0|auto_generated|mac_out4~DATAOUT3  = \Mult0|auto_generated|mac_out4_DATAOUT_bus [3];
assign \Mult0|auto_generated|mac_out4~DATAOUT4  = \Mult0|auto_generated|mac_out4_DATAOUT_bus [4];
assign \Mult0|auto_generated|mac_out4~DATAOUT5  = \Mult0|auto_generated|mac_out4_DATAOUT_bus [5];
assign \Mult0|auto_generated|mac_out4~DATAOUT6  = \Mult0|auto_generated|mac_out4_DATAOUT_bus [6];
assign \Mult0|auto_generated|mac_out4~DATAOUT7  = \Mult0|auto_generated|mac_out4_DATAOUT_bus [7];
assign \Mult0|auto_generated|mac_out4~DATAOUT8  = \Mult0|auto_generated|mac_out4_DATAOUT_bus [8];
assign \Mult0|auto_generated|mac_out4~DATAOUT9  = \Mult0|auto_generated|mac_out4_DATAOUT_bus [9];
assign \Mult0|auto_generated|mac_out4~DATAOUT10  = \Mult0|auto_generated|mac_out4_DATAOUT_bus [10];

assign \Mult0|auto_generated|mac_mult1~dataout  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [0];
assign \Mult0|auto_generated|mac_mult1~DATAOUT1  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [1];
assign \Mult0|auto_generated|mac_mult1~DATAOUT2  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [2];
assign \Mult0|auto_generated|mac_mult1~DATAOUT3  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [3];
assign \Mult0|auto_generated|mac_mult1~DATAOUT4  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [4];
assign \Mult0|auto_generated|mac_mult1~DATAOUT5  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [5];
assign \Mult0|auto_generated|mac_mult1~DATAOUT6  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [6];
assign \Mult0|auto_generated|mac_mult1~DATAOUT7  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [7];
assign \Mult0|auto_generated|mac_mult1~DATAOUT8  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [8];
assign \Mult0|auto_generated|mac_mult1~DATAOUT9  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [9];
assign \Mult0|auto_generated|mac_mult1~DATAOUT10  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [10];
assign \Mult0|auto_generated|mac_mult1~DATAOUT11  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [11];
assign \Mult0|auto_generated|mac_mult1~DATAOUT12  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [12];
assign \Mult0|auto_generated|mac_mult1~DATAOUT13  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [13];
assign \Mult0|auto_generated|mac_mult1~DATAOUT14  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [14];
assign \Mult0|auto_generated|mac_mult1~DATAOUT15  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [15];
assign \Mult0|auto_generated|mac_mult1~DATAOUT16  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [16];
assign \Mult0|auto_generated|mac_mult1~DATAOUT17  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [17];
assign \Mult0|auto_generated|mac_mult1~DATAOUT18  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [18];
assign \Mult0|auto_generated|mac_mult1~DATAOUT19  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [19];
assign \Mult0|auto_generated|mac_mult1~DATAOUT20  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [20];
assign \Mult0|auto_generated|mac_mult1~DATAOUT21  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [21];
assign \Mult0|auto_generated|mac_mult1~DATAOUT22  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [22];
assign \Mult0|auto_generated|mac_mult1~DATAOUT23  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [23];
assign \Mult0|auto_generated|mac_mult1~DATAOUT24  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [24];
assign \Mult0|auto_generated|mac_mult1~DATAOUT25  = \Mult0|auto_generated|mac_mult1_DATAOUT_bus [25];

assign \Mult0|auto_generated|mac_mult3~dataout  = \Mult0|auto_generated|mac_mult3_DATAOUT_bus [0];
assign \Mult0|auto_generated|mac_mult3~DATAOUT1  = \Mult0|auto_generated|mac_mult3_DATAOUT_bus [1];
assign \Mult0|auto_generated|mac_mult3~DATAOUT2  = \Mult0|auto_generated|mac_mult3_DATAOUT_bus [2];
assign \Mult0|auto_generated|mac_mult3~DATAOUT3  = \Mult0|auto_generated|mac_mult3_DATAOUT_bus [3];
assign \Mult0|auto_generated|mac_mult3~DATAOUT4  = \Mult0|auto_generated|mac_mult3_DATAOUT_bus [4];
assign \Mult0|auto_generated|mac_mult3~DATAOUT5  = \Mult0|auto_generated|mac_mult3_DATAOUT_bus [5];
assign \Mult0|auto_generated|mac_mult3~DATAOUT6  = \Mult0|auto_generated|mac_mult3_DATAOUT_bus [6];
assign \Mult0|auto_generated|mac_mult3~DATAOUT7  = \Mult0|auto_generated|mac_mult3_DATAOUT_bus [7];
assign \Mult0|auto_generated|mac_mult3~DATAOUT8  = \Mult0|auto_generated|mac_mult3_DATAOUT_bus [8];
assign \Mult0|auto_generated|mac_mult3~DATAOUT9  = \Mult0|auto_generated|mac_mult3_DATAOUT_bus [9];
assign \Mult0|auto_generated|mac_mult3~DATAOUT10  = \Mult0|auto_generated|mac_mult3_DATAOUT_bus [10];

lms_dsp_long_shift long_shift_inst(
	.q_b_0(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[0] ),
	.q_b_1(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[1] ),
	.q_b_2(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[2] ),
	.q_b_3(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[3] ),
	.q_b_4(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[4] ),
	.q_b_5(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[5] ),
	.q_b_6(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[6] ),
	.q_b_7(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[7] ),
	.q_b_8(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[8] ),
	.q_b_9(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[9] ),
	.q_b_10(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[10] ),
	.q_b_11(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[11] ),
	.q_b_12(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[12] ),
	.q_b_13(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[13] ),
	.q_b_14(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[14] ),
	.q_b_15(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[15] ),
	.q_b_01(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[0] ),
	.q_b_16(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[1] ),
	.q_b_21(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[2] ),
	.q_b_31(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[3] ),
	.q_b_41(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[4] ),
	.q_b_51(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[5] ),
	.q_b_61(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[6] ),
	.q_b_71(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[7] ),
	.q_b_81(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[8] ),
	.q_b_91(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[9] ),
	.q_b_101(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[10] ),
	.q_b_111(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[11] ),
	.q_b_121(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[12] ),
	.q_b_131(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[13] ),
	.q_b_141(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[14] ),
	.q_b_151(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[15] ),
	.always0(\always0~0_combout ),
	.delay_reg_24_0(delay_reg_24_0),
	.short_shift_full(\short_shift_full~q ),
	.short_to_long_arrived(\short_to_long_arrived~0_combout ),
	.GND_port(GND_port),
	.clk_clk(clk_clk));

lms_dsp_short_shift short_shift_inst(
	.mag_reg_0(mag_reg_0),
	.q_b_0(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[0] ),
	.mag_reg_1(mag_reg_1),
	.q_b_1(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[1] ),
	.mag_reg_2(mag_reg_2),
	.q_b_2(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[2] ),
	.mag_reg_3(mag_reg_3),
	.q_b_3(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[3] ),
	.mag_reg_4(mag_reg_4),
	.q_b_4(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[4] ),
	.mag_reg_5(mag_reg_5),
	.q_b_5(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[5] ),
	.mag_reg_6(mag_reg_6),
	.q_b_6(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[6] ),
	.mag_reg_7(mag_reg_7),
	.q_b_7(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[7] ),
	.mag_reg_8(mag_reg_8),
	.q_b_8(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[8] ),
	.mag_reg_9(mag_reg_9),
	.q_b_9(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[9] ),
	.mag_reg_10(mag_reg_10),
	.q_b_10(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[10] ),
	.mag_reg_11(mag_reg_11),
	.q_b_11(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[11] ),
	.mag_reg_12(mag_reg_12),
	.q_b_12(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[12] ),
	.q_b_13(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[13] ),
	.q_b_14(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[14] ),
	.q_b_15(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[15] ),
	.always0(\always0~2_combout ),
	.delay_reg_24_0(delay_reg_24_0),
	.GND_port(GND_port),
	.clk_clk(clk_clk));

dffeas \short_sum_reg[0] (
	.clk(clk_clk),
	.d(\short_sum_reg[0]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~2_combout ),
	.sload(gnd),
	.ena(\short_sum_reg[11]~20_combout ),
	.q(short_sum_reg_0),
	.prn(vcc));
defparam \short_sum_reg[0] .is_wysiwyg = "true";
defparam \short_sum_reg[0] .power_up = "low";

dffeas \short_sum_reg[1] (
	.clk(clk_clk),
	.d(\short_sum_reg[1]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~2_combout ),
	.sload(gnd),
	.ena(\short_sum_reg[11]~20_combout ),
	.q(short_sum_reg_1),
	.prn(vcc));
defparam \short_sum_reg[1] .is_wysiwyg = "true";
defparam \short_sum_reg[1] .power_up = "low";

dffeas \short_sum_reg[2] (
	.clk(clk_clk),
	.d(\short_sum_reg[2]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~2_combout ),
	.sload(gnd),
	.ena(\short_sum_reg[11]~20_combout ),
	.q(short_sum_reg_2),
	.prn(vcc));
defparam \short_sum_reg[2] .is_wysiwyg = "true";
defparam \short_sum_reg[2] .power_up = "low";

dffeas \short_sum_reg[3] (
	.clk(clk_clk),
	.d(\short_sum_reg[3]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~2_combout ),
	.sload(gnd),
	.ena(\short_sum_reg[11]~20_combout ),
	.q(short_sum_reg_3),
	.prn(vcc));
defparam \short_sum_reg[3] .is_wysiwyg = "true";
defparam \short_sum_reg[3] .power_up = "low";

dffeas \short_sum_reg[4] (
	.clk(clk_clk),
	.d(\short_sum_reg[4]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~2_combout ),
	.sload(gnd),
	.ena(\short_sum_reg[11]~20_combout ),
	.q(short_sum_reg_4),
	.prn(vcc));
defparam \short_sum_reg[4] .is_wysiwyg = "true";
defparam \short_sum_reg[4] .power_up = "low";

dffeas \short_sum_reg[5] (
	.clk(clk_clk),
	.d(\short_sum_reg[5]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~2_combout ),
	.sload(gnd),
	.ena(\short_sum_reg[11]~20_combout ),
	.q(short_sum_reg_5),
	.prn(vcc));
defparam \short_sum_reg[5] .is_wysiwyg = "true";
defparam \short_sum_reg[5] .power_up = "low";

dffeas \short_sum_reg[6] (
	.clk(clk_clk),
	.d(\short_sum_reg[6]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~2_combout ),
	.sload(gnd),
	.ena(\short_sum_reg[11]~20_combout ),
	.q(short_sum_reg_6),
	.prn(vcc));
defparam \short_sum_reg[6] .is_wysiwyg = "true";
defparam \short_sum_reg[6] .power_up = "low";

dffeas \short_sum_reg[7] (
	.clk(clk_clk),
	.d(\short_sum_reg[7]~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~2_combout ),
	.sload(gnd),
	.ena(\short_sum_reg[11]~20_combout ),
	.q(short_sum_reg_7),
	.prn(vcc));
defparam \short_sum_reg[7] .is_wysiwyg = "true";
defparam \short_sum_reg[7] .power_up = "low";

dffeas \short_sum_reg[8] (
	.clk(clk_clk),
	.d(\short_sum_reg[8]~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~2_combout ),
	.sload(gnd),
	.ena(\short_sum_reg[11]~20_combout ),
	.q(short_sum_reg_8),
	.prn(vcc));
defparam \short_sum_reg[8] .is_wysiwyg = "true";
defparam \short_sum_reg[8] .power_up = "low";

dffeas \short_sum_reg[9] (
	.clk(clk_clk),
	.d(\short_sum_reg[9]~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~2_combout ),
	.sload(gnd),
	.ena(\short_sum_reg[11]~20_combout ),
	.q(short_sum_reg_9),
	.prn(vcc));
defparam \short_sum_reg[9] .is_wysiwyg = "true";
defparam \short_sum_reg[9] .power_up = "low";

dffeas \short_sum_reg[10] (
	.clk(clk_clk),
	.d(\short_sum_reg[10]~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~2_combout ),
	.sload(gnd),
	.ena(\short_sum_reg[11]~20_combout ),
	.q(short_sum_reg_10),
	.prn(vcc));
defparam \short_sum_reg[10] .is_wysiwyg = "true";
defparam \short_sum_reg[10] .power_up = "low";

dffeas \short_sum_reg[11] (
	.clk(clk_clk),
	.d(\short_sum_reg[11]~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~2_combout ),
	.sload(gnd),
	.ena(\short_sum_reg[11]~20_combout ),
	.q(short_sum_reg_11),
	.prn(vcc));
defparam \short_sum_reg[11] .is_wysiwyg = "true";
defparam \short_sum_reg[11] .power_up = "low";

dffeas \short_sum_reg[12] (
	.clk(clk_clk),
	.d(\short_sum_reg[12]~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~2_combout ),
	.sload(gnd),
	.ena(\short_sum_reg[11]~20_combout ),
	.q(short_sum_reg_12),
	.prn(vcc));
defparam \short_sum_reg[12] .is_wysiwyg = "true";
defparam \short_sum_reg[12] .power_up = "low";

dffeas \short_sum_reg[13] (
	.clk(clk_clk),
	.d(\short_sum_reg[13]~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~2_combout ),
	.sload(gnd),
	.ena(\short_sum_reg[11]~20_combout ),
	.q(short_sum_reg_13),
	.prn(vcc));
defparam \short_sum_reg[13] .is_wysiwyg = "true";
defparam \short_sum_reg[13] .power_up = "low";

dffeas \short_sum_reg[14] (
	.clk(clk_clk),
	.d(\short_sum_reg[14]~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~2_combout ),
	.sload(gnd),
	.ena(\short_sum_reg[11]~20_combout ),
	.q(short_sum_reg_14),
	.prn(vcc));
defparam \short_sum_reg[14] .is_wysiwyg = "true";
defparam \short_sum_reg[14] .power_up = "low";

dffeas \short_sum_reg[15] (
	.clk(clk_clk),
	.d(\short_sum_reg[15]~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~2_combout ),
	.sload(gnd),
	.ena(\short_sum_reg[11]~20_combout ),
	.q(short_sum_reg_15),
	.prn(vcc));
defparam \short_sum_reg[15] .is_wysiwyg = "true";
defparam \short_sum_reg[15] .power_up = "low";

dffeas \short_sum_reg[16] (
	.clk(clk_clk),
	.d(\short_sum_reg[16]~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~2_combout ),
	.sload(gnd),
	.ena(\short_sum_reg[11]~20_combout ),
	.q(short_sum_reg_16),
	.prn(vcc));
defparam \short_sum_reg[16] .is_wysiwyg = "true";
defparam \short_sum_reg[16] .power_up = "low";

dffeas \short_sum_reg[17] (
	.clk(clk_clk),
	.d(\short_sum_reg[17]~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~2_combout ),
	.sload(gnd),
	.ena(\short_sum_reg[11]~20_combout ),
	.q(short_sum_reg_17),
	.prn(vcc));
defparam \short_sum_reg[17] .is_wysiwyg = "true";
defparam \short_sum_reg[17] .power_up = "low";

fiftyfivenm_lcell_comb \LessThan0~34 (
	.dataa(long_shift_rescale_17),
	.datab(short_sum_reg_17),
	.datac(gnd),
	.datad(gnd),
	.cin(\LessThan0~33_cout ),
	.combout(LessThan0),
	.cout());
defparam \LessThan0~34 .lut_mask = 16'hD4D4;
defparam \LessThan0~34 .sum_lutc_input = "cin";

dffeas \long_shift_rescale[0] (
	.clk(clk_clk),
	.d(\long_shift_rescale~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_0),
	.prn(vcc));
defparam \long_shift_rescale[0] .is_wysiwyg = "true";
defparam \long_shift_rescale[0] .power_up = "low";

dffeas \long_shift_rescale[1] (
	.clk(clk_clk),
	.d(\long_shift_rescale~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_1),
	.prn(vcc));
defparam \long_shift_rescale[1] .is_wysiwyg = "true";
defparam \long_shift_rescale[1] .power_up = "low";

dffeas \long_shift_rescale[2] (
	.clk(clk_clk),
	.d(\long_shift_rescale~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_2),
	.prn(vcc));
defparam \long_shift_rescale[2] .is_wysiwyg = "true";
defparam \long_shift_rescale[2] .power_up = "low";

dffeas \long_shift_rescale[3] (
	.clk(clk_clk),
	.d(\long_shift_rescale~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_3),
	.prn(vcc));
defparam \long_shift_rescale[3] .is_wysiwyg = "true";
defparam \long_shift_rescale[3] .power_up = "low";

dffeas \long_shift_rescale[4] (
	.clk(clk_clk),
	.d(\long_shift_rescale~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_4),
	.prn(vcc));
defparam \long_shift_rescale[4] .is_wysiwyg = "true";
defparam \long_shift_rescale[4] .power_up = "low";

dffeas \long_shift_rescale[5] (
	.clk(clk_clk),
	.d(\long_shift_rescale~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_5),
	.prn(vcc));
defparam \long_shift_rescale[5] .is_wysiwyg = "true";
defparam \long_shift_rescale[5] .power_up = "low";

dffeas \long_shift_rescale[6] (
	.clk(clk_clk),
	.d(\long_shift_rescale~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_6),
	.prn(vcc));
defparam \long_shift_rescale[6] .is_wysiwyg = "true";
defparam \long_shift_rescale[6] .power_up = "low";

dffeas \long_shift_rescale[7] (
	.clk(clk_clk),
	.d(\long_shift_rescale~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_7),
	.prn(vcc));
defparam \long_shift_rescale[7] .is_wysiwyg = "true";
defparam \long_shift_rescale[7] .power_up = "low";

dffeas \long_shift_rescale[8] (
	.clk(clk_clk),
	.d(\long_shift_rescale~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_8),
	.prn(vcc));
defparam \long_shift_rescale[8] .is_wysiwyg = "true";
defparam \long_shift_rescale[8] .power_up = "low";

dffeas \long_shift_rescale[9] (
	.clk(clk_clk),
	.d(\long_shift_rescale~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_9),
	.prn(vcc));
defparam \long_shift_rescale[9] .is_wysiwyg = "true";
defparam \long_shift_rescale[9] .power_up = "low";

dffeas \long_shift_rescale[10] (
	.clk(clk_clk),
	.d(\long_shift_rescale~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_10),
	.prn(vcc));
defparam \long_shift_rescale[10] .is_wysiwyg = "true";
defparam \long_shift_rescale[10] .power_up = "low";

dffeas \long_shift_rescale[11] (
	.clk(clk_clk),
	.d(\long_shift_rescale~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_11),
	.prn(vcc));
defparam \long_shift_rescale[11] .is_wysiwyg = "true";
defparam \long_shift_rescale[11] .power_up = "low";

dffeas \long_shift_rescale[12] (
	.clk(clk_clk),
	.d(\long_shift_rescale~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_12),
	.prn(vcc));
defparam \long_shift_rescale[12] .is_wysiwyg = "true";
defparam \long_shift_rescale[12] .power_up = "low";

dffeas \long_shift_rescale[13] (
	.clk(clk_clk),
	.d(\long_shift_rescale~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_13),
	.prn(vcc));
defparam \long_shift_rescale[13] .is_wysiwyg = "true";
defparam \long_shift_rescale[13] .power_up = "low";

dffeas \long_shift_rescale[14] (
	.clk(clk_clk),
	.d(\long_shift_rescale~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_14),
	.prn(vcc));
defparam \long_shift_rescale[14] .is_wysiwyg = "true";
defparam \long_shift_rescale[14] .power_up = "low";

dffeas \long_shift_rescale[15] (
	.clk(clk_clk),
	.d(\long_shift_rescale~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_15),
	.prn(vcc));
defparam \long_shift_rescale[15] .is_wysiwyg = "true";
defparam \long_shift_rescale[15] .power_up = "low";

dffeas \long_shift_rescale[16] (
	.clk(clk_clk),
	.d(\long_shift_rescale~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_16),
	.prn(vcc));
defparam \long_shift_rescale[16] .is_wysiwyg = "true";
defparam \long_shift_rescale[16] .power_up = "low";

dffeas \long_shift_rescale[17] (
	.clk(clk_clk),
	.d(\long_shift_rescale~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_17),
	.prn(vcc));
defparam \long_shift_rescale[17] .is_wysiwyg = "true";
defparam \long_shift_rescale[17] .power_up = "low";

dffeas \long_shift_rescale[18] (
	.clk(clk_clk),
	.d(\long_shift_rescale~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_18),
	.prn(vcc));
defparam \long_shift_rescale[18] .is_wysiwyg = "true";
defparam \long_shift_rescale[18] .power_up = "low";

dffeas \long_shift_rescale[19] (
	.clk(clk_clk),
	.d(\long_shift_rescale~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_19),
	.prn(vcc));
defparam \long_shift_rescale[19] .is_wysiwyg = "true";
defparam \long_shift_rescale[19] .power_up = "low";

dffeas \long_shift_rescale[20] (
	.clk(clk_clk),
	.d(\long_shift_rescale~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_20),
	.prn(vcc));
defparam \long_shift_rescale[20] .is_wysiwyg = "true";
defparam \long_shift_rescale[20] .power_up = "low";

fiftyfivenm_lcell_comb \launch~2 (
	.dataa(\Equal1~0_combout ),
	.datab(\Equal1~1_combout ),
	.datac(\launch~0_combout ),
	.datad(\launch~1_combout ),
	.cin(gnd),
	.combout(launch1),
	.cout());
defparam \launch~2 .lut_mask = 16'h8000;
defparam \launch~2 .sum_lutc_input = "datac";

dffeas \long_shift_rescale[25] (
	.clk(clk_clk),
	.d(\long_shift_rescale~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(long_shift_rescale_25),
	.prn(vcc));
defparam \long_shift_rescale[25] .is_wysiwyg = "true";
defparam \long_shift_rescale[25] .power_up = "low";

fiftyfivenm_lcell_comb launch(
	.dataa(LessThan0),
	.datab(launch1),
	.datac(gnd),
	.datad(long_shift_rescale_25),
	.cin(gnd),
	.combout(launch2),
	.cout());
defparam launch.lut_mask = 16'h0088;
defparam launch.sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~0 (
	.dataa(short_sum_reg_0),
	.datab(mag_reg_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
defparam \Add0~0 .lut_mask = 16'h6688;
defparam \Add0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \short_sum_reg[0]~18 (
	.dataa(\Add0~0_combout ),
	.datab(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[0] ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\short_sum_reg[0]~18_combout ),
	.cout(\short_sum_reg[0]~19 ));
defparam \short_sum_reg[0]~18 .lut_mask = 16'h66BB;
defparam \short_sum_reg[0]~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \always0~1 (
	.dataa(ppd_cfg_clear_rs),
	.datab(running_reg),
	.datac(gnd),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
defparam \always0~1 .lut_mask = 16'hEEFF;
defparam \always0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always0~2 (
	.dataa(\always0~1_combout ),
	.datab(LessThan0),
	.datac(launch1),
	.datad(long_shift_rescale_25),
	.cin(gnd),
	.combout(\always0~2_combout ),
	.cout());
defparam \always0~2 .lut_mask = 16'hAAEA;
defparam \always0~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \short_sum_reg[11]~20 (
	.dataa(\always0~2_combout ),
	.datab(delay_reg_24_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\short_sum_reg[11]~20_combout ),
	.cout());
defparam \short_sum_reg[11]~20 .lut_mask = 16'hEEEE;
defparam \short_sum_reg[11]~20 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~2 (
	.dataa(short_sum_reg_1),
	.datab(mag_reg_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'h9617;
defparam \Add0~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \short_sum_reg[1]~21 (
	.dataa(\Add0~2_combout ),
	.datab(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[1] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\short_sum_reg[0]~19 ),
	.combout(\short_sum_reg[1]~21_combout ),
	.cout(\short_sum_reg[1]~22 ));
defparam \short_sum_reg[1]~21 .lut_mask = 16'h694D;
defparam \short_sum_reg[1]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~4 (
	.dataa(short_sum_reg_2),
	.datab(mag_reg_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'h698E;
defparam \Add0~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \short_sum_reg[2]~23 (
	.dataa(\Add0~4_combout ),
	.datab(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[2] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\short_sum_reg[1]~22 ),
	.combout(\short_sum_reg[2]~23_combout ),
	.cout(\short_sum_reg[2]~24 ));
defparam \short_sum_reg[2]~23 .lut_mask = 16'h962B;
defparam \short_sum_reg[2]~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~6 (
	.dataa(short_sum_reg_3),
	.datab(mag_reg_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'h9617;
defparam \Add0~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \short_sum_reg[3]~25 (
	.dataa(\Add0~6_combout ),
	.datab(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[3] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\short_sum_reg[2]~24 ),
	.combout(\short_sum_reg[3]~25_combout ),
	.cout(\short_sum_reg[3]~26 ));
defparam \short_sum_reg[3]~25 .lut_mask = 16'h694D;
defparam \short_sum_reg[3]~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~8 (
	.dataa(short_sum_reg_4),
	.datab(mag_reg_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
defparam \Add0~8 .lut_mask = 16'h698E;
defparam \Add0~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \short_sum_reg[4]~27 (
	.dataa(\Add0~8_combout ),
	.datab(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[4] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\short_sum_reg[3]~26 ),
	.combout(\short_sum_reg[4]~27_combout ),
	.cout(\short_sum_reg[4]~28 ));
defparam \short_sum_reg[4]~27 .lut_mask = 16'h962B;
defparam \short_sum_reg[4]~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~10 (
	.dataa(short_sum_reg_5),
	.datab(mag_reg_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
defparam \Add0~10 .lut_mask = 16'h9617;
defparam \Add0~10 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \short_sum_reg[5]~29 (
	.dataa(\Add0~10_combout ),
	.datab(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[5] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\short_sum_reg[4]~28 ),
	.combout(\short_sum_reg[5]~29_combout ),
	.cout(\short_sum_reg[5]~30 ));
defparam \short_sum_reg[5]~29 .lut_mask = 16'h694D;
defparam \short_sum_reg[5]~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~12 (
	.dataa(short_sum_reg_6),
	.datab(mag_reg_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
defparam \Add0~12 .lut_mask = 16'h698E;
defparam \Add0~12 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \short_sum_reg[6]~31 (
	.dataa(\Add0~12_combout ),
	.datab(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[6] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\short_sum_reg[5]~30 ),
	.combout(\short_sum_reg[6]~31_combout ),
	.cout(\short_sum_reg[6]~32 ));
defparam \short_sum_reg[6]~31 .lut_mask = 16'h962B;
defparam \short_sum_reg[6]~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~14 (
	.dataa(short_sum_reg_7),
	.datab(mag_reg_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
defparam \Add0~14 .lut_mask = 16'h9617;
defparam \Add0~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \short_sum_reg[7]~33 (
	.dataa(\Add0~14_combout ),
	.datab(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[7] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\short_sum_reg[6]~32 ),
	.combout(\short_sum_reg[7]~33_combout ),
	.cout(\short_sum_reg[7]~34 ));
defparam \short_sum_reg[7]~33 .lut_mask = 16'h694D;
defparam \short_sum_reg[7]~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~16 (
	.dataa(short_sum_reg_8),
	.datab(mag_reg_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout(\Add0~17 ));
defparam \Add0~16 .lut_mask = 16'h698E;
defparam \Add0~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \short_sum_reg[8]~35 (
	.dataa(\Add0~16_combout ),
	.datab(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[8] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\short_sum_reg[7]~34 ),
	.combout(\short_sum_reg[8]~35_combout ),
	.cout(\short_sum_reg[8]~36 ));
defparam \short_sum_reg[8]~35 .lut_mask = 16'h962B;
defparam \short_sum_reg[8]~35 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~18 (
	.dataa(short_sum_reg_9),
	.datab(mag_reg_9),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~17 ),
	.combout(\Add0~18_combout ),
	.cout(\Add0~19 ));
defparam \Add0~18 .lut_mask = 16'h9617;
defparam \Add0~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \short_sum_reg[9]~37 (
	.dataa(\Add0~18_combout ),
	.datab(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[9] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\short_sum_reg[8]~36 ),
	.combout(\short_sum_reg[9]~37_combout ),
	.cout(\short_sum_reg[9]~38 ));
defparam \short_sum_reg[9]~37 .lut_mask = 16'h694D;
defparam \short_sum_reg[9]~37 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~20 (
	.dataa(short_sum_reg_10),
	.datab(mag_reg_10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~19 ),
	.combout(\Add0~20_combout ),
	.cout(\Add0~21 ));
defparam \Add0~20 .lut_mask = 16'h698E;
defparam \Add0~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \short_sum_reg[10]~39 (
	.dataa(\Add0~20_combout ),
	.datab(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[10] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\short_sum_reg[9]~38 ),
	.combout(\short_sum_reg[10]~39_combout ),
	.cout(\short_sum_reg[10]~40 ));
defparam \short_sum_reg[10]~39 .lut_mask = 16'h962B;
defparam \short_sum_reg[10]~39 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~22 (
	.dataa(short_sum_reg_11),
	.datab(mag_reg_11),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~21 ),
	.combout(\Add0~22_combout ),
	.cout(\Add0~23 ));
defparam \Add0~22 .lut_mask = 16'h9617;
defparam \Add0~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \short_sum_reg[11]~41 (
	.dataa(\Add0~22_combout ),
	.datab(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[11] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\short_sum_reg[10]~40 ),
	.combout(\short_sum_reg[11]~41_combout ),
	.cout(\short_sum_reg[11]~42 ));
defparam \short_sum_reg[11]~41 .lut_mask = 16'h694D;
defparam \short_sum_reg[11]~41 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~24 (
	.dataa(short_sum_reg_12),
	.datab(mag_reg_12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~23 ),
	.combout(\Add0~24_combout ),
	.cout(\Add0~25 ));
defparam \Add0~24 .lut_mask = 16'h698E;
defparam \Add0~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \short_sum_reg[12]~43 (
	.dataa(\Add0~24_combout ),
	.datab(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[12] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\short_sum_reg[11]~42 ),
	.combout(\short_sum_reg[12]~43_combout ),
	.cout(\short_sum_reg[12]~44 ));
defparam \short_sum_reg[12]~43 .lut_mask = 16'h962B;
defparam \short_sum_reg[12]~43 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~26 (
	.dataa(short_sum_reg_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~25 ),
	.combout(\Add0~26_combout ),
	.cout(\Add0~27 ));
defparam \Add0~26 .lut_mask = 16'h5A5F;
defparam \Add0~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \short_sum_reg[13]~45 (
	.dataa(\Add0~26_combout ),
	.datab(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[13] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\short_sum_reg[12]~44 ),
	.combout(\short_sum_reg[13]~45_combout ),
	.cout(\short_sum_reg[13]~46 ));
defparam \short_sum_reg[13]~45 .lut_mask = 16'h694D;
defparam \short_sum_reg[13]~45 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~28 (
	.dataa(short_sum_reg_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~27 ),
	.combout(\Add0~28_combout ),
	.cout(\Add0~29 ));
defparam \Add0~28 .lut_mask = 16'hA50A;
defparam \Add0~28 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \short_sum_reg[14]~47 (
	.dataa(\Add0~28_combout ),
	.datab(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[14] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\short_sum_reg[13]~46 ),
	.combout(\short_sum_reg[14]~47_combout ),
	.cout(\short_sum_reg[14]~48 ));
defparam \short_sum_reg[14]~47 .lut_mask = 16'h962B;
defparam \short_sum_reg[14]~47 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~30 (
	.dataa(short_sum_reg_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~29 ),
	.combout(\Add0~30_combout ),
	.cout(\Add0~31 ));
defparam \Add0~30 .lut_mask = 16'h5A5F;
defparam \Add0~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \short_sum_reg[15]~49 (
	.dataa(\Add0~30_combout ),
	.datab(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[15] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\short_sum_reg[14]~48 ),
	.combout(\short_sum_reg[15]~49_combout ),
	.cout(\short_sum_reg[15]~50 ));
defparam \short_sum_reg[15]~49 .lut_mask = 16'h694D;
defparam \short_sum_reg[15]~49 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~32 (
	.dataa(short_sum_reg_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~31 ),
	.combout(\Add0~32_combout ),
	.cout(\Add0~33 ));
defparam \Add0~32 .lut_mask = 16'hA50A;
defparam \Add0~32 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \short_sum_reg[16]~51 (
	.dataa(\Add0~32_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\short_sum_reg[15]~50 ),
	.combout(\short_sum_reg[16]~51_combout ),
	.cout(\short_sum_reg[16]~52 ));
defparam \short_sum_reg[16]~51 .lut_mask = 16'h5AAF;
defparam \short_sum_reg[16]~51 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~34 (
	.dataa(short_sum_reg_17),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~33 ),
	.combout(\Add0~34_combout ),
	.cout());
defparam \Add0~34 .lut_mask = 16'h5A5A;
defparam \Add0~34 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \short_sum_reg[17]~53 (
	.dataa(\Add0~34_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\short_sum_reg[16]~52 ),
	.combout(\short_sum_reg[17]~53_combout ),
	.cout());
defparam \short_sum_reg[17]~53 .lut_mask = 16'hA5A5;
defparam \short_sum_reg[17]~53 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~1 (
	.dataa(long_shift_rescale_0),
	.datab(short_sum_reg_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan0~1_cout ));
defparam \LessThan0~1 .lut_mask = 16'h0044;
defparam \LessThan0~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~3 (
	.dataa(long_shift_rescale_1),
	.datab(short_sum_reg_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~1_cout ),
	.combout(),
	.cout(\LessThan0~3_cout ));
defparam \LessThan0~3 .lut_mask = 16'h002B;
defparam \LessThan0~3 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~5 (
	.dataa(long_shift_rescale_2),
	.datab(short_sum_reg_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~3_cout ),
	.combout(),
	.cout(\LessThan0~5_cout ));
defparam \LessThan0~5 .lut_mask = 16'h004D;
defparam \LessThan0~5 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~7 (
	.dataa(long_shift_rescale_3),
	.datab(short_sum_reg_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~5_cout ),
	.combout(),
	.cout(\LessThan0~7_cout ));
defparam \LessThan0~7 .lut_mask = 16'h002B;
defparam \LessThan0~7 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~9 (
	.dataa(long_shift_rescale_4),
	.datab(short_sum_reg_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~7_cout ),
	.combout(),
	.cout(\LessThan0~9_cout ));
defparam \LessThan0~9 .lut_mask = 16'h004D;
defparam \LessThan0~9 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~11 (
	.dataa(long_shift_rescale_5),
	.datab(short_sum_reg_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~9_cout ),
	.combout(),
	.cout(\LessThan0~11_cout ));
defparam \LessThan0~11 .lut_mask = 16'h002B;
defparam \LessThan0~11 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~13 (
	.dataa(long_shift_rescale_6),
	.datab(short_sum_reg_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~11_cout ),
	.combout(),
	.cout(\LessThan0~13_cout ));
defparam \LessThan0~13 .lut_mask = 16'h004D;
defparam \LessThan0~13 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~15 (
	.dataa(long_shift_rescale_7),
	.datab(short_sum_reg_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~13_cout ),
	.combout(),
	.cout(\LessThan0~15_cout ));
defparam \LessThan0~15 .lut_mask = 16'h002B;
defparam \LessThan0~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~17 (
	.dataa(long_shift_rescale_8),
	.datab(short_sum_reg_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~15_cout ),
	.combout(),
	.cout(\LessThan0~17_cout ));
defparam \LessThan0~17 .lut_mask = 16'h004D;
defparam \LessThan0~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~19 (
	.dataa(long_shift_rescale_9),
	.datab(short_sum_reg_9),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~17_cout ),
	.combout(),
	.cout(\LessThan0~19_cout ));
defparam \LessThan0~19 .lut_mask = 16'h002B;
defparam \LessThan0~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~21 (
	.dataa(long_shift_rescale_10),
	.datab(short_sum_reg_10),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~19_cout ),
	.combout(),
	.cout(\LessThan0~21_cout ));
defparam \LessThan0~21 .lut_mask = 16'h004D;
defparam \LessThan0~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~23 (
	.dataa(long_shift_rescale_11),
	.datab(short_sum_reg_11),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~21_cout ),
	.combout(),
	.cout(\LessThan0~23_cout ));
defparam \LessThan0~23 .lut_mask = 16'h002B;
defparam \LessThan0~23 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~25 (
	.dataa(long_shift_rescale_12),
	.datab(short_sum_reg_12),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~23_cout ),
	.combout(),
	.cout(\LessThan0~25_cout ));
defparam \LessThan0~25 .lut_mask = 16'h004D;
defparam \LessThan0~25 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~27 (
	.dataa(long_shift_rescale_13),
	.datab(short_sum_reg_13),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~25_cout ),
	.combout(),
	.cout(\LessThan0~27_cout ));
defparam \LessThan0~27 .lut_mask = 16'h002B;
defparam \LessThan0~27 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~29 (
	.dataa(long_shift_rescale_14),
	.datab(short_sum_reg_14),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~27_cout ),
	.combout(),
	.cout(\LessThan0~29_cout ));
defparam \LessThan0~29 .lut_mask = 16'h004D;
defparam \LessThan0~29 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~31 (
	.dataa(long_shift_rescale_15),
	.datab(short_sum_reg_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~29_cout ),
	.combout(),
	.cout(\LessThan0~31_cout ));
defparam \LessThan0~31 .lut_mask = 16'h002B;
defparam \LessThan0~31 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~33 (
	.dataa(long_shift_rescale_16),
	.datab(short_sum_reg_16),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~31_cout ),
	.combout(),
	.cout(\LessThan0~33_cout ));
defparam \LessThan0~33 .lut_mask = 16'h004D;
defparam \LessThan0~33 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add3~0 (
	.dataa(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[0] ),
	.datab(\long_sum_reg[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add3~0_combout ),
	.cout(\Add3~1 ));
defparam \Add3~0 .lut_mask = 16'h6688;
defparam \Add3~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \long_sum_reg[0]~21 (
	.dataa(\Add3~0_combout ),
	.datab(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[0] ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\long_sum_reg[0]~21_combout ),
	.cout(\long_sum_reg[0]~22 ));
defparam \long_sum_reg[0]~21 .lut_mask = 16'h66BB;
defparam \long_sum_reg[0]~21 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \always0~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(gnd),
	.datac(gnd),
	.datad(ppd_cfg_clear_rs),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hFF55;
defparam \always0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \short_counter[0]~5 (
	.dataa(\short_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\short_counter[0]~5_combout ),
	.cout(\short_counter[0]~6 ));
defparam \short_counter[0]~5 .lut_mask = 16'h55AA;
defparam \short_counter[0]~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \short_to_long_arrived~0 (
	.dataa(delay_reg_24_0),
	.datab(\short_shift_full~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\short_to_long_arrived~0_combout ),
	.cout());
defparam \short_to_long_arrived~0 .lut_mask = 16'h8888;
defparam \short_to_long_arrived~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \short_to_long_arrived~1 (
	.dataa(\short_to_long_arrived~q ),
	.datab(\short_to_long_arrived~0_combout ),
	.datac(\Equal0~1_combout ),
	.datad(\always0~2_combout ),
	.cin(gnd),
	.combout(\short_to_long_arrived~1_combout ),
	.cout());
defparam \short_to_long_arrived~1 .lut_mask = 16'h00EA;
defparam \short_to_long_arrived~1 .sum_lutc_input = "datac";

dffeas short_to_long_arrived(
	.clk(clk_clk),
	.d(\short_to_long_arrived~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\short_to_long_arrived~q ),
	.prn(vcc));
defparam short_to_long_arrived.is_wysiwyg = "true";
defparam short_to_long_arrived.power_up = "low";

fiftyfivenm_lcell_comb \short_counter[0]~15 (
	.dataa(\short_to_long_arrived~q ),
	.datab(\always0~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\short_counter[0]~15_combout ),
	.cout());
defparam \short_counter[0]~15 .lut_mask = 16'hEEEE;
defparam \short_counter[0]~15 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \short_counter[0]~16 (
	.dataa(\short_to_long_arrived~q ),
	.datab(\short_shift_full~q ),
	.datac(\Equal0~1_combout ),
	.datad(delay_reg_24_0),
	.cin(gnd),
	.combout(\short_counter[0]~16_combout ),
	.cout());
defparam \short_counter[0]~16 .lut_mask = 16'h8AFF;
defparam \short_counter[0]~16 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \short_counter[0]~17 (
	.dataa(\short_counter[0]~16_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\always0~2_combout ),
	.cin(gnd),
	.combout(\short_counter[0]~17_combout ),
	.cout());
defparam \short_counter[0]~17 .lut_mask = 16'hFF55;
defparam \short_counter[0]~17 .sum_lutc_input = "datac";

dffeas \short_counter[0] (
	.clk(clk_clk),
	.d(\short_counter[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\short_counter[0]~15_combout ),
	.sload(gnd),
	.ena(\short_counter[0]~17_combout ),
	.q(\short_counter[0]~q ),
	.prn(vcc));
defparam \short_counter[0] .is_wysiwyg = "true";
defparam \short_counter[0] .power_up = "low";

fiftyfivenm_lcell_comb \short_counter[1]~7 (
	.dataa(\short_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\short_counter[0]~6 ),
	.combout(\short_counter[1]~7_combout ),
	.cout(\short_counter[1]~8 ));
defparam \short_counter[1]~7 .lut_mask = 16'h5A5F;
defparam \short_counter[1]~7 .sum_lutc_input = "cin";

dffeas \short_counter[1] (
	.clk(clk_clk),
	.d(\short_counter[1]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\short_counter[0]~15_combout ),
	.sload(gnd),
	.ena(\short_counter[0]~17_combout ),
	.q(\short_counter[1]~q ),
	.prn(vcc));
defparam \short_counter[1] .is_wysiwyg = "true";
defparam \short_counter[1] .power_up = "low";

fiftyfivenm_lcell_comb \short_counter[2]~9 (
	.dataa(\short_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\short_counter[1]~8 ),
	.combout(\short_counter[2]~9_combout ),
	.cout(\short_counter[2]~10 ));
defparam \short_counter[2]~9 .lut_mask = 16'hA50A;
defparam \short_counter[2]~9 .sum_lutc_input = "cin";

dffeas \short_counter[2] (
	.clk(clk_clk),
	.d(\short_counter[2]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\short_counter[0]~15_combout ),
	.sload(gnd),
	.ena(\short_counter[0]~17_combout ),
	.q(\short_counter[2]~q ),
	.prn(vcc));
defparam \short_counter[2] .is_wysiwyg = "true";
defparam \short_counter[2] .power_up = "low";

fiftyfivenm_lcell_comb \short_counter[3]~11 (
	.dataa(\short_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\short_counter[2]~10 ),
	.combout(\short_counter[3]~11_combout ),
	.cout(\short_counter[3]~12 ));
defparam \short_counter[3]~11 .lut_mask = 16'h5A5F;
defparam \short_counter[3]~11 .sum_lutc_input = "cin";

dffeas \short_counter[3] (
	.clk(clk_clk),
	.d(\short_counter[3]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\short_counter[0]~15_combout ),
	.sload(gnd),
	.ena(\short_counter[0]~17_combout ),
	.q(\short_counter[3]~q ),
	.prn(vcc));
defparam \short_counter[3] .is_wysiwyg = "true";
defparam \short_counter[3] .power_up = "low";

fiftyfivenm_lcell_comb \short_counter[4]~13 (
	.dataa(\short_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\short_counter[3]~12 ),
	.combout(\short_counter[4]~13_combout ),
	.cout());
defparam \short_counter[4]~13 .lut_mask = 16'hA5A5;
defparam \short_counter[4]~13 .sum_lutc_input = "cin";

dffeas \short_counter[4] (
	.clk(clk_clk),
	.d(\short_counter[4]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\short_counter[0]~15_combout ),
	.sload(gnd),
	.ena(\short_counter[0]~17_combout ),
	.q(\short_counter[4]~q ),
	.prn(vcc));
defparam \short_counter[4] .is_wysiwyg = "true";
defparam \short_counter[4] .power_up = "low";

fiftyfivenm_lcell_comb \Equal0~0 (
	.dataa(\short_counter[0]~q ),
	.datab(\short_counter[1]~q ),
	.datac(\short_counter[2]~q ),
	.datad(\short_counter[3]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h8000;
defparam \Equal0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal0~1 (
	.dataa(\short_counter[4]~q ),
	.datab(\Equal0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h8888;
defparam \Equal0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \short_shift_full~0 (
	.dataa(\short_shift_full~q ),
	.datab(delay_reg_24_0),
	.datac(\Equal0~1_combout ),
	.datad(\always0~2_combout ),
	.cin(gnd),
	.combout(\short_shift_full~0_combout ),
	.cout());
defparam \short_shift_full~0 .lut_mask = 16'h00EA;
defparam \short_shift_full~0 .sum_lutc_input = "datac";

dffeas short_shift_full(
	.clk(clk_clk),
	.d(\short_shift_full~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\short_shift_full~q ),
	.prn(vcc));
defparam short_shift_full.is_wysiwyg = "true";
defparam short_shift_full.power_up = "low";

fiftyfivenm_lcell_comb \long_sum_reg[1]~23 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(delay_reg_24_0),
	.datac(\short_shift_full~q ),
	.datad(ppd_cfg_clear_rs),
	.cin(gnd),
	.combout(\long_sum_reg[1]~23_combout ),
	.cout());
defparam \long_sum_reg[1]~23 .lut_mask = 16'hFFD5;
defparam \long_sum_reg[1]~23 .sum_lutc_input = "datac";

dffeas \long_sum_reg[0] (
	.clk(clk_clk),
	.d(\long_sum_reg[0]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[0]~q ),
	.prn(vcc));
defparam \long_sum_reg[0] .is_wysiwyg = "true";
defparam \long_sum_reg[0] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~2 (
	.dataa(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[1] ),
	.datab(\long_sum_reg[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~1 ),
	.combout(\Add3~2_combout ),
	.cout(\Add3~3 ));
defparam \Add3~2 .lut_mask = 16'h9617;
defparam \Add3~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[1]~24 (
	.dataa(\Add3~2_combout ),
	.datab(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[1] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_sum_reg[0]~22 ),
	.combout(\long_sum_reg[1]~24_combout ),
	.cout(\long_sum_reg[1]~25 ));
defparam \long_sum_reg[1]~24 .lut_mask = 16'h694D;
defparam \long_sum_reg[1]~24 .sum_lutc_input = "cin";

dffeas \long_sum_reg[1] (
	.clk(clk_clk),
	.d(\long_sum_reg[1]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[1]~q ),
	.prn(vcc));
defparam \long_sum_reg[1] .is_wysiwyg = "true";
defparam \long_sum_reg[1] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~4 (
	.dataa(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[2] ),
	.datab(\long_sum_reg[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~3 ),
	.combout(\Add3~4_combout ),
	.cout(\Add3~5 ));
defparam \Add3~4 .lut_mask = 16'h698E;
defparam \Add3~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[2]~26 (
	.dataa(\Add3~4_combout ),
	.datab(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[2] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_sum_reg[1]~25 ),
	.combout(\long_sum_reg[2]~26_combout ),
	.cout(\long_sum_reg[2]~27 ));
defparam \long_sum_reg[2]~26 .lut_mask = 16'h962B;
defparam \long_sum_reg[2]~26 .sum_lutc_input = "cin";

dffeas \long_sum_reg[2] (
	.clk(clk_clk),
	.d(\long_sum_reg[2]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[2]~q ),
	.prn(vcc));
defparam \long_sum_reg[2] .is_wysiwyg = "true";
defparam \long_sum_reg[2] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~6 (
	.dataa(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[3] ),
	.datab(\long_sum_reg[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~5 ),
	.combout(\Add3~6_combout ),
	.cout(\Add3~7 ));
defparam \Add3~6 .lut_mask = 16'h9617;
defparam \Add3~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[3]~28 (
	.dataa(\Add3~6_combout ),
	.datab(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[3] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_sum_reg[2]~27 ),
	.combout(\long_sum_reg[3]~28_combout ),
	.cout(\long_sum_reg[3]~29 ));
defparam \long_sum_reg[3]~28 .lut_mask = 16'h694D;
defparam \long_sum_reg[3]~28 .sum_lutc_input = "cin";

dffeas \long_sum_reg[3] (
	.clk(clk_clk),
	.d(\long_sum_reg[3]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[3]~q ),
	.prn(vcc));
defparam \long_sum_reg[3] .is_wysiwyg = "true";
defparam \long_sum_reg[3] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~8 (
	.dataa(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[4] ),
	.datab(\long_sum_reg[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~7 ),
	.combout(\Add3~8_combout ),
	.cout(\Add3~9 ));
defparam \Add3~8 .lut_mask = 16'h698E;
defparam \Add3~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[4]~30 (
	.dataa(\Add3~8_combout ),
	.datab(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[4] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_sum_reg[3]~29 ),
	.combout(\long_sum_reg[4]~30_combout ),
	.cout(\long_sum_reg[4]~31 ));
defparam \long_sum_reg[4]~30 .lut_mask = 16'h962B;
defparam \long_sum_reg[4]~30 .sum_lutc_input = "cin";

dffeas \long_sum_reg[4] (
	.clk(clk_clk),
	.d(\long_sum_reg[4]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[4]~q ),
	.prn(vcc));
defparam \long_sum_reg[4] .is_wysiwyg = "true";
defparam \long_sum_reg[4] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~10 (
	.dataa(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[5] ),
	.datab(\long_sum_reg[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~9 ),
	.combout(\Add3~10_combout ),
	.cout(\Add3~11 ));
defparam \Add3~10 .lut_mask = 16'h9617;
defparam \Add3~10 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[5]~32 (
	.dataa(\Add3~10_combout ),
	.datab(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[5] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_sum_reg[4]~31 ),
	.combout(\long_sum_reg[5]~32_combout ),
	.cout(\long_sum_reg[5]~33 ));
defparam \long_sum_reg[5]~32 .lut_mask = 16'h694D;
defparam \long_sum_reg[5]~32 .sum_lutc_input = "cin";

dffeas \long_sum_reg[5] (
	.clk(clk_clk),
	.d(\long_sum_reg[5]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[5]~q ),
	.prn(vcc));
defparam \long_sum_reg[5] .is_wysiwyg = "true";
defparam \long_sum_reg[5] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~12 (
	.dataa(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[6] ),
	.datab(\long_sum_reg[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~11 ),
	.combout(\Add3~12_combout ),
	.cout(\Add3~13 ));
defparam \Add3~12 .lut_mask = 16'h698E;
defparam \Add3~12 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[6]~34 (
	.dataa(\Add3~12_combout ),
	.datab(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[6] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_sum_reg[5]~33 ),
	.combout(\long_sum_reg[6]~34_combout ),
	.cout(\long_sum_reg[6]~35 ));
defparam \long_sum_reg[6]~34 .lut_mask = 16'h962B;
defparam \long_sum_reg[6]~34 .sum_lutc_input = "cin";

dffeas \long_sum_reg[6] (
	.clk(clk_clk),
	.d(\long_sum_reg[6]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[6]~q ),
	.prn(vcc));
defparam \long_sum_reg[6] .is_wysiwyg = "true";
defparam \long_sum_reg[6] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~14 (
	.dataa(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[7] ),
	.datab(\long_sum_reg[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~13 ),
	.combout(\Add3~14_combout ),
	.cout(\Add3~15 ));
defparam \Add3~14 .lut_mask = 16'h9617;
defparam \Add3~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[7]~36 (
	.dataa(\Add3~14_combout ),
	.datab(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[7] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_sum_reg[6]~35 ),
	.combout(\long_sum_reg[7]~36_combout ),
	.cout(\long_sum_reg[7]~37 ));
defparam \long_sum_reg[7]~36 .lut_mask = 16'h694D;
defparam \long_sum_reg[7]~36 .sum_lutc_input = "cin";

dffeas \long_sum_reg[7] (
	.clk(clk_clk),
	.d(\long_sum_reg[7]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[7]~q ),
	.prn(vcc));
defparam \long_sum_reg[7] .is_wysiwyg = "true";
defparam \long_sum_reg[7] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~16 (
	.dataa(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[8] ),
	.datab(\long_sum_reg[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~15 ),
	.combout(\Add3~16_combout ),
	.cout(\Add3~17 ));
defparam \Add3~16 .lut_mask = 16'h698E;
defparam \Add3~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[8]~38 (
	.dataa(\Add3~16_combout ),
	.datab(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[8] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_sum_reg[7]~37 ),
	.combout(\long_sum_reg[8]~38_combout ),
	.cout(\long_sum_reg[8]~39 ));
defparam \long_sum_reg[8]~38 .lut_mask = 16'h962B;
defparam \long_sum_reg[8]~38 .sum_lutc_input = "cin";

dffeas \long_sum_reg[8] (
	.clk(clk_clk),
	.d(\long_sum_reg[8]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[8]~q ),
	.prn(vcc));
defparam \long_sum_reg[8] .is_wysiwyg = "true";
defparam \long_sum_reg[8] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~18 (
	.dataa(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[9] ),
	.datab(\long_sum_reg[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~17 ),
	.combout(\Add3~18_combout ),
	.cout(\Add3~19 ));
defparam \Add3~18 .lut_mask = 16'h9617;
defparam \Add3~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[9]~40 (
	.dataa(\Add3~18_combout ),
	.datab(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[9] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_sum_reg[8]~39 ),
	.combout(\long_sum_reg[9]~40_combout ),
	.cout(\long_sum_reg[9]~41 ));
defparam \long_sum_reg[9]~40 .lut_mask = 16'h694D;
defparam \long_sum_reg[9]~40 .sum_lutc_input = "cin";

dffeas \long_sum_reg[9] (
	.clk(clk_clk),
	.d(\long_sum_reg[9]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[9]~q ),
	.prn(vcc));
defparam \long_sum_reg[9] .is_wysiwyg = "true";
defparam \long_sum_reg[9] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~20 (
	.dataa(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[10] ),
	.datab(\long_sum_reg[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~19 ),
	.combout(\Add3~20_combout ),
	.cout(\Add3~21 ));
defparam \Add3~20 .lut_mask = 16'h698E;
defparam \Add3~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[10]~42 (
	.dataa(\Add3~20_combout ),
	.datab(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[10] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_sum_reg[9]~41 ),
	.combout(\long_sum_reg[10]~42_combout ),
	.cout(\long_sum_reg[10]~43 ));
defparam \long_sum_reg[10]~42 .lut_mask = 16'h962B;
defparam \long_sum_reg[10]~42 .sum_lutc_input = "cin";

dffeas \long_sum_reg[10] (
	.clk(clk_clk),
	.d(\long_sum_reg[10]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[10]~q ),
	.prn(vcc));
defparam \long_sum_reg[10] .is_wysiwyg = "true";
defparam \long_sum_reg[10] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~22 (
	.dataa(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[11] ),
	.datab(\long_sum_reg[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~21 ),
	.combout(\Add3~22_combout ),
	.cout(\Add3~23 ));
defparam \Add3~22 .lut_mask = 16'h9617;
defparam \Add3~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[11]~44 (
	.dataa(\Add3~22_combout ),
	.datab(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[11] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_sum_reg[10]~43 ),
	.combout(\long_sum_reg[11]~44_combout ),
	.cout(\long_sum_reg[11]~45 ));
defparam \long_sum_reg[11]~44 .lut_mask = 16'h694D;
defparam \long_sum_reg[11]~44 .sum_lutc_input = "cin";

dffeas \long_sum_reg[11] (
	.clk(clk_clk),
	.d(\long_sum_reg[11]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[11]~q ),
	.prn(vcc));
defparam \long_sum_reg[11] .is_wysiwyg = "true";
defparam \long_sum_reg[11] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~24 (
	.dataa(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[12] ),
	.datab(\long_sum_reg[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~23 ),
	.combout(\Add3~24_combout ),
	.cout(\Add3~25 ));
defparam \Add3~24 .lut_mask = 16'h698E;
defparam \Add3~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[12]~46 (
	.dataa(\Add3~24_combout ),
	.datab(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[12] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_sum_reg[11]~45 ),
	.combout(\long_sum_reg[12]~46_combout ),
	.cout(\long_sum_reg[12]~47 ));
defparam \long_sum_reg[12]~46 .lut_mask = 16'h962B;
defparam \long_sum_reg[12]~46 .sum_lutc_input = "cin";

dffeas \long_sum_reg[12] (
	.clk(clk_clk),
	.d(\long_sum_reg[12]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[12]~q ),
	.prn(vcc));
defparam \long_sum_reg[12] .is_wysiwyg = "true";
defparam \long_sum_reg[12] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~26 (
	.dataa(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[13] ),
	.datab(\long_sum_reg[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~25 ),
	.combout(\Add3~26_combout ),
	.cout(\Add3~27 ));
defparam \Add3~26 .lut_mask = 16'h9617;
defparam \Add3~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[13]~48 (
	.dataa(\Add3~26_combout ),
	.datab(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[13] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_sum_reg[12]~47 ),
	.combout(\long_sum_reg[13]~48_combout ),
	.cout(\long_sum_reg[13]~49 ));
defparam \long_sum_reg[13]~48 .lut_mask = 16'h694D;
defparam \long_sum_reg[13]~48 .sum_lutc_input = "cin";

dffeas \long_sum_reg[13] (
	.clk(clk_clk),
	.d(\long_sum_reg[13]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[13]~q ),
	.prn(vcc));
defparam \long_sum_reg[13] .is_wysiwyg = "true";
defparam \long_sum_reg[13] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~28 (
	.dataa(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[14] ),
	.datab(\long_sum_reg[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~27 ),
	.combout(\Add3~28_combout ),
	.cout(\Add3~29 ));
defparam \Add3~28 .lut_mask = 16'h698E;
defparam \Add3~28 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[14]~50 (
	.dataa(\Add3~28_combout ),
	.datab(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[14] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_sum_reg[13]~49 ),
	.combout(\long_sum_reg[14]~50_combout ),
	.cout(\long_sum_reg[14]~51 ));
defparam \long_sum_reg[14]~50 .lut_mask = 16'h962B;
defparam \long_sum_reg[14]~50 .sum_lutc_input = "cin";

dffeas \long_sum_reg[14] (
	.clk(clk_clk),
	.d(\long_sum_reg[14]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[14]~q ),
	.prn(vcc));
defparam \long_sum_reg[14] .is_wysiwyg = "true";
defparam \long_sum_reg[14] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~30 (
	.dataa(\short_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[15] ),
	.datab(\long_sum_reg[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~29 ),
	.combout(\Add3~30_combout ),
	.cout(\Add3~31 ));
defparam \Add3~30 .lut_mask = 16'h9617;
defparam \Add3~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[15]~52 (
	.dataa(\Add3~30_combout ),
	.datab(\long_shift_inst|ALTSHIFT_TAPS_component|auto_generated|altsyncram2|q_b[15] ),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_sum_reg[14]~51 ),
	.combout(\long_sum_reg[15]~52_combout ),
	.cout(\long_sum_reg[15]~53 ));
defparam \long_sum_reg[15]~52 .lut_mask = 16'h694D;
defparam \long_sum_reg[15]~52 .sum_lutc_input = "cin";

dffeas \long_sum_reg[15] (
	.clk(clk_clk),
	.d(\long_sum_reg[15]~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[15]~q ),
	.prn(vcc));
defparam \long_sum_reg[15] .is_wysiwyg = "true";
defparam \long_sum_reg[15] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~32 (
	.dataa(\long_sum_reg[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~31 ),
	.combout(\Add3~32_combout ),
	.cout(\Add3~33 ));
defparam \Add3~32 .lut_mask = 16'hA50A;
defparam \Add3~32 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[16]~54 (
	.dataa(\Add3~32_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_sum_reg[15]~53 ),
	.combout(\long_sum_reg[16]~54_combout ),
	.cout(\long_sum_reg[16]~55 ));
defparam \long_sum_reg[16]~54 .lut_mask = 16'h5AAF;
defparam \long_sum_reg[16]~54 .sum_lutc_input = "cin";

dffeas \long_sum_reg[16] (
	.clk(clk_clk),
	.d(\long_sum_reg[16]~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[16]~q ),
	.prn(vcc));
defparam \long_sum_reg[16] .is_wysiwyg = "true";
defparam \long_sum_reg[16] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~34 (
	.dataa(\long_sum_reg[17]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~33 ),
	.combout(\Add3~34_combout ),
	.cout(\Add3~35 ));
defparam \Add3~34 .lut_mask = 16'h5A5F;
defparam \Add3~34 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[17]~56 (
	.dataa(\Add3~34_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_sum_reg[16]~55 ),
	.combout(\long_sum_reg[17]~56_combout ),
	.cout(\long_sum_reg[17]~57 ));
defparam \long_sum_reg[17]~56 .lut_mask = 16'hA505;
defparam \long_sum_reg[17]~56 .sum_lutc_input = "cin";

dffeas \long_sum_reg[17] (
	.clk(clk_clk),
	.d(\long_sum_reg[17]~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[17]~q ),
	.prn(vcc));
defparam \long_sum_reg[17] .is_wysiwyg = "true";
defparam \long_sum_reg[17] .power_up = "low";

fiftyfivenm_mac_mult \Mult0|auto_generated|mac_mult1 (
	.signa(gnd),
	.signb(gnd),
	.clk(gnd),
	.aclr(gnd),
	.ena(vcc),
	.dataa({\long_sum_reg[17]~q ,\long_sum_reg[16]~q ,\long_sum_reg[15]~q ,\long_sum_reg[14]~q ,\long_sum_reg[13]~q ,\long_sum_reg[12]~q ,\long_sum_reg[11]~q ,\long_sum_reg[10]~q ,\long_sum_reg[9]~q ,\long_sum_reg[8]~q ,\long_sum_reg[7]~q ,\long_sum_reg[6]~q ,\long_sum_reg[5]~q ,
\long_sum_reg[4]~q ,\long_sum_reg[3]~q ,\long_sum_reg[2]~q ,\long_sum_reg[1]~q ,\long_sum_reg[0]~q }),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ppd_cfg_threshold_7,ppd_cfg_threshold_6,ppd_cfg_threshold_5,ppd_cfg_threshold_4,ppd_cfg_threshold_3,ppd_cfg_threshold_2,ppd_cfg_threshold_1,ppd_cfg_threshold_0}),
	.dataout(\Mult0|auto_generated|mac_mult1_DATAOUT_bus ));
defparam \Mult0|auto_generated|mac_mult1 .dataa_clock = "none";
defparam \Mult0|auto_generated|mac_mult1 .dataa_width = 18;
defparam \Mult0|auto_generated|mac_mult1 .datab_clock = "none";
defparam \Mult0|auto_generated|mac_mult1 .datab_width = 8;
defparam \Mult0|auto_generated|mac_mult1 .signa_clock = "none";
defparam \Mult0|auto_generated|mac_mult1 .signb_clock = "none";

fiftyfivenm_mac_out \Mult0|auto_generated|mac_out2 (
	.clk(gnd),
	.aclr(gnd),
	.ena(vcc),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Mult0|auto_generated|mac_mult1~DATAOUT25 ,\Mult0|auto_generated|mac_mult1~DATAOUT24 ,\Mult0|auto_generated|mac_mult1~DATAOUT23 ,\Mult0|auto_generated|mac_mult1~DATAOUT22 ,\Mult0|auto_generated|mac_mult1~DATAOUT21 ,
\Mult0|auto_generated|mac_mult1~DATAOUT20 ,\Mult0|auto_generated|mac_mult1~DATAOUT19 ,\Mult0|auto_generated|mac_mult1~DATAOUT18 ,\Mult0|auto_generated|mac_mult1~DATAOUT17 ,\Mult0|auto_generated|mac_mult1~DATAOUT16 ,\Mult0|auto_generated|mac_mult1~DATAOUT15 ,
\Mult0|auto_generated|mac_mult1~DATAOUT14 ,\Mult0|auto_generated|mac_mult1~DATAOUT13 ,\Mult0|auto_generated|mac_mult1~DATAOUT12 ,\Mult0|auto_generated|mac_mult1~DATAOUT11 ,\Mult0|auto_generated|mac_mult1~DATAOUT10 ,\Mult0|auto_generated|mac_mult1~DATAOUT9 ,
\Mult0|auto_generated|mac_mult1~DATAOUT8 ,\Mult0|auto_generated|mac_mult1~DATAOUT7 ,\Mult0|auto_generated|mac_mult1~DATAOUT6 ,\Mult0|auto_generated|mac_mult1~DATAOUT5 ,\Mult0|auto_generated|mac_mult1~DATAOUT4 ,\Mult0|auto_generated|mac_mult1~DATAOUT3 ,
\Mult0|auto_generated|mac_mult1~DATAOUT2 ,\Mult0|auto_generated|mac_mult1~DATAOUT1 ,\Mult0|auto_generated|mac_mult1~dataout }),
	.dataout(\Mult0|auto_generated|mac_out2_DATAOUT_bus ));
defparam \Mult0|auto_generated|mac_out2 .dataa_width = 26;
defparam \Mult0|auto_generated|mac_out2 .output_clock = "none";

fiftyfivenm_lcell_comb \long_shift_rescale~22 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Mult0|auto_generated|w138w[3] ),
	.datac(gnd),
	.datad(ppd_cfg_clear_rs),
	.cin(gnd),
	.combout(\long_shift_rescale~22_combout ),
	.cout());
defparam \long_shift_rescale~22 .lut_mask = 16'h0088;
defparam \long_shift_rescale~22 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \long_shift_rescale~23 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Mult0|auto_generated|w138w[4] ),
	.datac(gnd),
	.datad(ppd_cfg_clear_rs),
	.cin(gnd),
	.combout(\long_shift_rescale~23_combout ),
	.cout());
defparam \long_shift_rescale~23 .lut_mask = 16'h0088;
defparam \long_shift_rescale~23 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \long_shift_rescale~24 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Mult0|auto_generated|w138w[5] ),
	.datac(gnd),
	.datad(ppd_cfg_clear_rs),
	.cin(gnd),
	.combout(\long_shift_rescale~24_combout ),
	.cout());
defparam \long_shift_rescale~24 .lut_mask = 16'h0088;
defparam \long_shift_rescale~24 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \long_shift_rescale~25 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Mult0|auto_generated|w138w[6] ),
	.datac(gnd),
	.datad(ppd_cfg_clear_rs),
	.cin(gnd),
	.combout(\long_shift_rescale~25_combout ),
	.cout());
defparam \long_shift_rescale~25 .lut_mask = 16'h0088;
defparam \long_shift_rescale~25 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \long_shift_rescale~26 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Mult0|auto_generated|w138w[7] ),
	.datac(gnd),
	.datad(ppd_cfg_clear_rs),
	.cin(gnd),
	.combout(\long_shift_rescale~26_combout ),
	.cout());
defparam \long_shift_rescale~26 .lut_mask = 16'h0088;
defparam \long_shift_rescale~26 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \long_shift_rescale~27 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Mult0|auto_generated|w138w[8] ),
	.datac(gnd),
	.datad(ppd_cfg_clear_rs),
	.cin(gnd),
	.combout(\long_shift_rescale~27_combout ),
	.cout());
defparam \long_shift_rescale~27 .lut_mask = 16'h0088;
defparam \long_shift_rescale~27 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \long_shift_rescale~28 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Mult0|auto_generated|w138w[9] ),
	.datac(gnd),
	.datad(ppd_cfg_clear_rs),
	.cin(gnd),
	.combout(\long_shift_rescale~28_combout ),
	.cout());
defparam \long_shift_rescale~28 .lut_mask = 16'h0088;
defparam \long_shift_rescale~28 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \long_shift_rescale~29 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Mult0|auto_generated|w138w[10] ),
	.datac(gnd),
	.datad(ppd_cfg_clear_rs),
	.cin(gnd),
	.combout(\long_shift_rescale~29_combout ),
	.cout());
defparam \long_shift_rescale~29 .lut_mask = 16'h0088;
defparam \long_shift_rescale~29 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \long_shift_rescale~30 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Mult0|auto_generated|w138w[11] ),
	.datac(gnd),
	.datad(ppd_cfg_clear_rs),
	.cin(gnd),
	.combout(\long_shift_rescale~30_combout ),
	.cout());
defparam \long_shift_rescale~30 .lut_mask = 16'h0088;
defparam \long_shift_rescale~30 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \long_shift_rescale~31 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Mult0|auto_generated|w138w[12] ),
	.datac(gnd),
	.datad(ppd_cfg_clear_rs),
	.cin(gnd),
	.combout(\long_shift_rescale~31_combout ),
	.cout());
defparam \long_shift_rescale~31 .lut_mask = 16'h0088;
defparam \long_shift_rescale~31 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \long_shift_rescale~32 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Mult0|auto_generated|w138w[13] ),
	.datac(gnd),
	.datad(ppd_cfg_clear_rs),
	.cin(gnd),
	.combout(\long_shift_rescale~32_combout ),
	.cout());
defparam \long_shift_rescale~32 .lut_mask = 16'h0088;
defparam \long_shift_rescale~32 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \long_shift_rescale~33 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Mult0|auto_generated|w138w[14] ),
	.datac(gnd),
	.datad(ppd_cfg_clear_rs),
	.cin(gnd),
	.combout(\long_shift_rescale~33_combout ),
	.cout());
defparam \long_shift_rescale~33 .lut_mask = 16'h0088;
defparam \long_shift_rescale~33 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \long_shift_rescale~34 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Mult0|auto_generated|w138w[15] ),
	.datac(gnd),
	.datad(ppd_cfg_clear_rs),
	.cin(gnd),
	.combout(\long_shift_rescale~34_combout ),
	.cout());
defparam \long_shift_rescale~34 .lut_mask = 16'h0088;
defparam \long_shift_rescale~34 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \long_shift_rescale~35 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Mult0|auto_generated|w138w[16] ),
	.datac(gnd),
	.datad(ppd_cfg_clear_rs),
	.cin(gnd),
	.combout(\long_shift_rescale~35_combout ),
	.cout());
defparam \long_shift_rescale~35 .lut_mask = 16'h0088;
defparam \long_shift_rescale~35 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \long_shift_rescale~36 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Mult0|auto_generated|w138w[17] ),
	.datac(gnd),
	.datad(ppd_cfg_clear_rs),
	.cin(gnd),
	.combout(\long_shift_rescale~36_combout ),
	.cout());
defparam \long_shift_rescale~36 .lut_mask = 16'h0088;
defparam \long_shift_rescale~36 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add3~36 (
	.dataa(\long_sum_reg[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~35 ),
	.combout(\Add3~36_combout ),
	.cout(\Add3~37 ));
defparam \Add3~36 .lut_mask = 16'hA50A;
defparam \Add3~36 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[18]~58 (
	.dataa(\Add3~36_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_sum_reg[17]~57 ),
	.combout(\long_sum_reg[18]~58_combout ),
	.cout(\long_sum_reg[18]~59 ));
defparam \long_sum_reg[18]~58 .lut_mask = 16'h5AAF;
defparam \long_sum_reg[18]~58 .sum_lutc_input = "cin";

dffeas \long_sum_reg[18] (
	.clk(clk_clk),
	.d(\long_sum_reg[18]~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[18]~q ),
	.prn(vcc));
defparam \long_sum_reg[18] .is_wysiwyg = "true";
defparam \long_sum_reg[18] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~38 (
	.dataa(\long_sum_reg[19]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~37 ),
	.combout(\Add3~38_combout ),
	.cout(\Add3~39 ));
defparam \Add3~38 .lut_mask = 16'h5A5F;
defparam \Add3~38 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[19]~60 (
	.dataa(\Add3~38_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_sum_reg[18]~59 ),
	.combout(\long_sum_reg[19]~60_combout ),
	.cout(\long_sum_reg[19]~61 ));
defparam \long_sum_reg[19]~60 .lut_mask = 16'hA505;
defparam \long_sum_reg[19]~60 .sum_lutc_input = "cin";

dffeas \long_sum_reg[19] (
	.clk(clk_clk),
	.d(\long_sum_reg[19]~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[19]~q ),
	.prn(vcc));
defparam \long_sum_reg[19] .is_wysiwyg = "true";
defparam \long_sum_reg[19] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~40 (
	.dataa(\long_sum_reg[20]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add3~39 ),
	.combout(\Add3~40_combout ),
	.cout());
defparam \Add3~40 .lut_mask = 16'hA5A5;
defparam \Add3~40 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_sum_reg[20]~62 (
	.dataa(\Add3~40_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\long_sum_reg[19]~61 ),
	.combout(\long_sum_reg[20]~62_combout ),
	.cout());
defparam \long_sum_reg[20]~62 .lut_mask = 16'h5A5A;
defparam \long_sum_reg[20]~62 .sum_lutc_input = "cin";

dffeas \long_sum_reg[20] (
	.clk(clk_clk),
	.d(\long_sum_reg[20]~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_sum_reg[1]~23_combout ),
	.q(\long_sum_reg[20]~q ),
	.prn(vcc));
defparam \long_sum_reg[20] .is_wysiwyg = "true";
defparam \long_sum_reg[20] .power_up = "low";

fiftyfivenm_mac_mult \Mult0|auto_generated|mac_mult3 (
	.signa(gnd),
	.signb(gnd),
	.clk(gnd),
	.aclr(gnd),
	.ena(vcc),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\long_sum_reg[20]~q ,\long_sum_reg[19]~q ,\long_sum_reg[18]~q }),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ppd_cfg_threshold_7,ppd_cfg_threshold_6,ppd_cfg_threshold_5,ppd_cfg_threshold_4,ppd_cfg_threshold_3,ppd_cfg_threshold_2,ppd_cfg_threshold_1,ppd_cfg_threshold_0}),
	.dataout(\Mult0|auto_generated|mac_mult3_DATAOUT_bus ));
defparam \Mult0|auto_generated|mac_mult3 .dataa_clock = "none";
defparam \Mult0|auto_generated|mac_mult3 .dataa_width = 3;
defparam \Mult0|auto_generated|mac_mult3 .datab_clock = "none";
defparam \Mult0|auto_generated|mac_mult3 .datab_width = 8;
defparam \Mult0|auto_generated|mac_mult3 .signa_clock = "none";
defparam \Mult0|auto_generated|mac_mult3 .signb_clock = "none";

fiftyfivenm_mac_out \Mult0|auto_generated|mac_out4 (
	.clk(gnd),
	.aclr(gnd),
	.ena(vcc),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Mult0|auto_generated|mac_mult3~DATAOUT10 ,\Mult0|auto_generated|mac_mult3~DATAOUT9 ,\Mult0|auto_generated|mac_mult3~DATAOUT8 ,\Mult0|auto_generated|mac_mult3~DATAOUT7 ,
\Mult0|auto_generated|mac_mult3~DATAOUT6 ,\Mult0|auto_generated|mac_mult3~DATAOUT5 ,\Mult0|auto_generated|mac_mult3~DATAOUT4 ,\Mult0|auto_generated|mac_mult3~DATAOUT3 ,\Mult0|auto_generated|mac_mult3~DATAOUT2 ,\Mult0|auto_generated|mac_mult3~DATAOUT1 ,
\Mult0|auto_generated|mac_mult3~dataout }),
	.dataout(\Mult0|auto_generated|mac_out4_DATAOUT_bus ));
defparam \Mult0|auto_generated|mac_out4 .dataa_width = 11;
defparam \Mult0|auto_generated|mac_out4 .output_clock = "none";

fiftyfivenm_lcell_comb \Mult0|auto_generated|op_1~0 (
	.dataa(\Mult0|auto_generated|mac_out4~dataout ),
	.datab(\Mult0|auto_generated|mac_out2~DATAOUT18 ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Mult0|auto_generated|op_1~0_combout ),
	.cout(\Mult0|auto_generated|op_1~1 ));
defparam \Mult0|auto_generated|op_1~0 .lut_mask = 16'h6688;
defparam \Mult0|auto_generated|op_1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \long_shift_rescale~37 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(ppd_cfg_clear_rs),
	.datac(\Mult0|auto_generated|op_1~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\long_shift_rescale~37_combout ),
	.cout());
defparam \long_shift_rescale~37 .lut_mask = 16'h2020;
defparam \long_shift_rescale~37 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mult0|auto_generated|op_1~2 (
	.dataa(\Mult0|auto_generated|mac_out4~DATAOUT1 ),
	.datab(\Mult0|auto_generated|mac_out2~DATAOUT19 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mult0|auto_generated|op_1~1 ),
	.combout(\Mult0|auto_generated|op_1~2_combout ),
	.cout(\Mult0|auto_generated|op_1~3 ));
defparam \Mult0|auto_generated|op_1~2 .lut_mask = 16'h9617;
defparam \Mult0|auto_generated|op_1~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_shift_rescale~38 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(ppd_cfg_clear_rs),
	.datac(\Mult0|auto_generated|op_1~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\long_shift_rescale~38_combout ),
	.cout());
defparam \long_shift_rescale~38 .lut_mask = 16'h2020;
defparam \long_shift_rescale~38 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mult0|auto_generated|op_1~4 (
	.dataa(\Mult0|auto_generated|mac_out4~DATAOUT2 ),
	.datab(\Mult0|auto_generated|mac_out2~DATAOUT20 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mult0|auto_generated|op_1~3 ),
	.combout(\Mult0|auto_generated|op_1~4_combout ),
	.cout(\Mult0|auto_generated|op_1~5 ));
defparam \Mult0|auto_generated|op_1~4 .lut_mask = 16'h698E;
defparam \Mult0|auto_generated|op_1~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_shift_rescale~39 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(ppd_cfg_clear_rs),
	.datac(\Mult0|auto_generated|op_1~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\long_shift_rescale~39_combout ),
	.cout());
defparam \long_shift_rescale~39 .lut_mask = 16'h2020;
defparam \long_shift_rescale~39 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mult0|auto_generated|op_1~6 (
	.dataa(\Mult0|auto_generated|mac_out4~DATAOUT3 ),
	.datab(\Mult0|auto_generated|mac_out2~DATAOUT21 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mult0|auto_generated|op_1~5 ),
	.combout(\Mult0|auto_generated|op_1~6_combout ),
	.cout(\Mult0|auto_generated|op_1~7 ));
defparam \Mult0|auto_generated|op_1~6 .lut_mask = 16'h9617;
defparam \Mult0|auto_generated|op_1~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_shift_rescale~40 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(ppd_cfg_clear_rs),
	.datac(\Mult0|auto_generated|op_1~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\long_shift_rescale~40_combout ),
	.cout());
defparam \long_shift_rescale~40 .lut_mask = 16'h2020;
defparam \long_shift_rescale~40 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mult0|auto_generated|op_1~8 (
	.dataa(\Mult0|auto_generated|mac_out4~DATAOUT4 ),
	.datab(\Mult0|auto_generated|mac_out2~DATAOUT22 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mult0|auto_generated|op_1~7 ),
	.combout(\Mult0|auto_generated|op_1~8_combout ),
	.cout(\Mult0|auto_generated|op_1~9 ));
defparam \Mult0|auto_generated|op_1~8 .lut_mask = 16'h698E;
defparam \Mult0|auto_generated|op_1~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_shift_rescale~41 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(ppd_cfg_clear_rs),
	.datac(\Mult0|auto_generated|op_1~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\long_shift_rescale~41_combout ),
	.cout());
defparam \long_shift_rescale~41 .lut_mask = 16'h2020;
defparam \long_shift_rescale~41 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mult0|auto_generated|op_1~10 (
	.dataa(\Mult0|auto_generated|mac_out4~DATAOUT5 ),
	.datab(\Mult0|auto_generated|mac_out2~DATAOUT23 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mult0|auto_generated|op_1~9 ),
	.combout(\Mult0|auto_generated|op_1~10_combout ),
	.cout(\Mult0|auto_generated|op_1~11 ));
defparam \Mult0|auto_generated|op_1~10 .lut_mask = 16'h9617;
defparam \Mult0|auto_generated|op_1~10 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_shift_rescale~42 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(ppd_cfg_clear_rs),
	.datac(\Mult0|auto_generated|op_1~10_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\long_shift_rescale~42_combout ),
	.cout());
defparam \long_shift_rescale~42 .lut_mask = 16'h2020;
defparam \long_shift_rescale~42 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \long_counter[0]~8 (
	.dataa(\long_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\long_counter[0]~8_combout ),
	.cout(\long_counter[0]~9 ));
defparam \long_counter[0]~8 .lut_mask = 16'h55AA;
defparam \long_counter[0]~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \long_counter[1]~11 (
	.dataa(\long_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_counter[0]~9 ),
	.combout(\long_counter[1]~11_combout ),
	.cout(\long_counter[1]~12 ));
defparam \long_counter[1]~11 .lut_mask = 16'h5A5F;
defparam \long_counter[1]~11 .sum_lutc_input = "cin";

dffeas \long_counter[1] (
	.clk(clk_clk),
	.d(\long_counter[1]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_counter[0]~10_combout ),
	.q(\long_counter[1]~q ),
	.prn(vcc));
defparam \long_counter[1] .is_wysiwyg = "true";
defparam \long_counter[1] .power_up = "low";

fiftyfivenm_lcell_comb \long_counter[2]~13 (
	.dataa(\long_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_counter[1]~12 ),
	.combout(\long_counter[2]~13_combout ),
	.cout(\long_counter[2]~14 ));
defparam \long_counter[2]~13 .lut_mask = 16'hA50A;
defparam \long_counter[2]~13 .sum_lutc_input = "cin";

dffeas \long_counter[2] (
	.clk(clk_clk),
	.d(\long_counter[2]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_counter[0]~10_combout ),
	.q(\long_counter[2]~q ),
	.prn(vcc));
defparam \long_counter[2] .is_wysiwyg = "true";
defparam \long_counter[2] .power_up = "low";

fiftyfivenm_lcell_comb \long_counter[3]~15 (
	.dataa(\long_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_counter[2]~14 ),
	.combout(\long_counter[3]~15_combout ),
	.cout(\long_counter[3]~16 ));
defparam \long_counter[3]~15 .lut_mask = 16'h5A5F;
defparam \long_counter[3]~15 .sum_lutc_input = "cin";

dffeas \long_counter[3] (
	.clk(clk_clk),
	.d(\long_counter[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_counter[0]~10_combout ),
	.q(\long_counter[3]~q ),
	.prn(vcc));
defparam \long_counter[3] .is_wysiwyg = "true";
defparam \long_counter[3] .power_up = "low";

fiftyfivenm_lcell_comb \long_counter[4]~17 (
	.dataa(\long_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_counter[3]~16 ),
	.combout(\long_counter[4]~17_combout ),
	.cout(\long_counter[4]~18 ));
defparam \long_counter[4]~17 .lut_mask = 16'hA50A;
defparam \long_counter[4]~17 .sum_lutc_input = "cin";

dffeas \long_counter[4] (
	.clk(clk_clk),
	.d(\long_counter[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_counter[0]~10_combout ),
	.q(\long_counter[4]~q ),
	.prn(vcc));
defparam \long_counter[4] .is_wysiwyg = "true";
defparam \long_counter[4] .power_up = "low";

fiftyfivenm_lcell_comb \long_counter[5]~19 (
	.dataa(\long_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_counter[4]~18 ),
	.combout(\long_counter[5]~19_combout ),
	.cout(\long_counter[5]~20 ));
defparam \long_counter[5]~19 .lut_mask = 16'h5A5F;
defparam \long_counter[5]~19 .sum_lutc_input = "cin";

dffeas \long_counter[5] (
	.clk(clk_clk),
	.d(\long_counter[5]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_counter[0]~10_combout ),
	.q(\long_counter[5]~q ),
	.prn(vcc));
defparam \long_counter[5] .is_wysiwyg = "true";
defparam \long_counter[5] .power_up = "low";

fiftyfivenm_lcell_comb \long_counter[6]~21 (
	.dataa(\long_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\long_counter[5]~20 ),
	.combout(\long_counter[6]~21_combout ),
	.cout(\long_counter[6]~22 ));
defparam \long_counter[6]~21 .lut_mask = 16'hA50A;
defparam \long_counter[6]~21 .sum_lutc_input = "cin";

dffeas \long_counter[6] (
	.clk(clk_clk),
	.d(\long_counter[6]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_counter[0]~10_combout ),
	.q(\long_counter[6]~q ),
	.prn(vcc));
defparam \long_counter[6] .is_wysiwyg = "true";
defparam \long_counter[6] .power_up = "low";

fiftyfivenm_lcell_comb \long_counter[7]~23 (
	.dataa(\long_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\long_counter[6]~22 ),
	.combout(\long_counter[7]~23_combout ),
	.cout());
defparam \long_counter[7]~23 .lut_mask = 16'h5A5A;
defparam \long_counter[7]~23 .sum_lutc_input = "cin";

dffeas \long_counter[7] (
	.clk(clk_clk),
	.d(\long_counter[7]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_counter[0]~10_combout ),
	.q(\long_counter[7]~q ),
	.prn(vcc));
defparam \long_counter[7] .is_wysiwyg = "true";
defparam \long_counter[7] .power_up = "low";

fiftyfivenm_lcell_comb \Equal1~1 (
	.dataa(\long_counter[4]~q ),
	.datab(\long_counter[5]~q ),
	.datac(\long_counter[6]~q ),
	.datad(\long_counter[7]~q ),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
defparam \Equal1~1 .lut_mask = 16'h8000;
defparam \Equal1~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \long_counter[0]~10 (
	.dataa(\always0~0_combout ),
	.datab(\Equal1~0_combout ),
	.datac(\Equal1~1_combout ),
	.datad(\short_to_long_arrived~0_combout ),
	.cin(gnd),
	.combout(\long_counter[0]~10_combout ),
	.cout());
defparam \long_counter[0]~10 .lut_mask = 16'hBFAA;
defparam \long_counter[0]~10 .sum_lutc_input = "datac";

dffeas \long_counter[0] (
	.clk(clk_clk),
	.d(\long_counter[0]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always0~0_combout ),
	.sload(gnd),
	.ena(\long_counter[0]~10_combout ),
	.q(\long_counter[0]~q ),
	.prn(vcc));
defparam \long_counter[0] .is_wysiwyg = "true";
defparam \long_counter[0] .power_up = "low";

fiftyfivenm_lcell_comb \Equal1~0 (
	.dataa(\long_counter[0]~q ),
	.datab(\long_counter[1]~q ),
	.datac(\long_counter[2]~q ),
	.datad(\long_counter[3]~q ),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'h8000;
defparam \Equal1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \launch~0 (
	.dataa(\short_to_long_arrived~q ),
	.datab(long_shift_rescale_18),
	.datac(long_shift_rescale_19),
	.datad(long_shift_rescale_20),
	.cin(gnd),
	.combout(\launch~0_combout ),
	.cout());
defparam \launch~0 .lut_mask = 16'h0002;
defparam \launch~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mult0|auto_generated|op_1~12 (
	.dataa(\Mult0|auto_generated|mac_out4~DATAOUT6 ),
	.datab(\Mult0|auto_generated|mac_out2~DATAOUT24 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mult0|auto_generated|op_1~11 ),
	.combout(\Mult0|auto_generated|op_1~12_combout ),
	.cout(\Mult0|auto_generated|op_1~13 ));
defparam \Mult0|auto_generated|op_1~12 .lut_mask = 16'h698E;
defparam \Mult0|auto_generated|op_1~12 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_shift_rescale~43 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(ppd_cfg_clear_rs),
	.datac(\Mult0|auto_generated|op_1~12_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\long_shift_rescale~43_combout ),
	.cout());
defparam \long_shift_rescale~43 .lut_mask = 16'h2020;
defparam \long_shift_rescale~43 .sum_lutc_input = "datac";

dffeas \long_shift_rescale[21] (
	.clk(clk_clk),
	.d(\long_shift_rescale~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\long_shift_rescale[21]~q ),
	.prn(vcc));
defparam \long_shift_rescale[21] .is_wysiwyg = "true";
defparam \long_shift_rescale[21] .power_up = "low";

fiftyfivenm_lcell_comb \Mult0|auto_generated|op_1~14 (
	.dataa(\Mult0|auto_generated|mac_out4~DATAOUT7 ),
	.datab(\Mult0|auto_generated|mac_out2~DATAOUT25 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mult0|auto_generated|op_1~13 ),
	.combout(\Mult0|auto_generated|op_1~14_combout ),
	.cout(\Mult0|auto_generated|op_1~15 ));
defparam \Mult0|auto_generated|op_1~14 .lut_mask = 16'h9617;
defparam \Mult0|auto_generated|op_1~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_shift_rescale~44 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(ppd_cfg_clear_rs),
	.datac(\Mult0|auto_generated|op_1~14_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\long_shift_rescale~44_combout ),
	.cout());
defparam \long_shift_rescale~44 .lut_mask = 16'h2020;
defparam \long_shift_rescale~44 .sum_lutc_input = "datac";

dffeas \long_shift_rescale[22] (
	.clk(clk_clk),
	.d(\long_shift_rescale~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\long_shift_rescale[22]~q ),
	.prn(vcc));
defparam \long_shift_rescale[22] .is_wysiwyg = "true";
defparam \long_shift_rescale[22] .power_up = "low";

fiftyfivenm_lcell_comb \Mult0|auto_generated|op_1~16 (
	.dataa(\Mult0|auto_generated|mac_out4~DATAOUT8 ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mult0|auto_generated|op_1~15 ),
	.combout(\Mult0|auto_generated|op_1~16_combout ),
	.cout(\Mult0|auto_generated|op_1~17 ));
defparam \Mult0|auto_generated|op_1~16 .lut_mask = 16'hA50A;
defparam \Mult0|auto_generated|op_1~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_shift_rescale~45 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(ppd_cfg_clear_rs),
	.datac(\Mult0|auto_generated|op_1~16_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\long_shift_rescale~45_combout ),
	.cout());
defparam \long_shift_rescale~45 .lut_mask = 16'h2020;
defparam \long_shift_rescale~45 .sum_lutc_input = "datac";

dffeas \long_shift_rescale[23] (
	.clk(clk_clk),
	.d(\long_shift_rescale~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\long_shift_rescale[23]~q ),
	.prn(vcc));
defparam \long_shift_rescale[23] .is_wysiwyg = "true";
defparam \long_shift_rescale[23] .power_up = "low";

fiftyfivenm_lcell_comb \Mult0|auto_generated|op_1~18 (
	.dataa(\Mult0|auto_generated|mac_out4~DATAOUT9 ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mult0|auto_generated|op_1~17 ),
	.combout(\Mult0|auto_generated|op_1~18_combout ),
	.cout(\Mult0|auto_generated|op_1~19 ));
defparam \Mult0|auto_generated|op_1~18 .lut_mask = 16'h5A5F;
defparam \Mult0|auto_generated|op_1~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_shift_rescale~46 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(ppd_cfg_clear_rs),
	.datac(\Mult0|auto_generated|op_1~18_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\long_shift_rescale~46_combout ),
	.cout());
defparam \long_shift_rescale~46 .lut_mask = 16'h2020;
defparam \long_shift_rescale~46 .sum_lutc_input = "datac";

dffeas \long_shift_rescale[24] (
	.clk(clk_clk),
	.d(\long_shift_rescale~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\long_shift_rescale[24]~q ),
	.prn(vcc));
defparam \long_shift_rescale[24] .is_wysiwyg = "true";
defparam \long_shift_rescale[24] .power_up = "low";

fiftyfivenm_lcell_comb \launch~1 (
	.dataa(\long_shift_rescale[21]~q ),
	.datab(\long_shift_rescale[22]~q ),
	.datac(\long_shift_rescale[23]~q ),
	.datad(\long_shift_rescale[24]~q ),
	.cin(gnd),
	.combout(\launch~1_combout ),
	.cout());
defparam \launch~1 .lut_mask = 16'h0001;
defparam \launch~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mult0|auto_generated|op_1~20 (
	.dataa(\Mult0|auto_generated|mac_out4~DATAOUT10 ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Mult0|auto_generated|op_1~19 ),
	.combout(\Mult0|auto_generated|op_1~20_combout ),
	.cout());
defparam \Mult0|auto_generated|op_1~20 .lut_mask = 16'hA5A5;
defparam \Mult0|auto_generated|op_1~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \long_shift_rescale~47 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(ppd_cfg_clear_rs),
	.datac(\Mult0|auto_generated|op_1~20_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\long_shift_rescale~47_combout ),
	.cout());
defparam \long_shift_rescale~47 .lut_mask = 16'h2020;
defparam \long_shift_rescale~47 .sum_lutc_input = "datac";

endmodule

module lms_dsp_long_shift (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_01,
	q_b_16,
	q_b_21,
	q_b_31,
	q_b_41,
	q_b_51,
	q_b_61,
	q_b_71,
	q_b_81,
	q_b_91,
	q_b_101,
	q_b_111,
	q_b_121,
	q_b_131,
	q_b_141,
	q_b_151,
	always0,
	delay_reg_24_0,
	short_shift_full,
	short_to_long_arrived,
	GND_port,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	q_b_0;
input 	q_b_1;
input 	q_b_2;
input 	q_b_3;
input 	q_b_4;
input 	q_b_5;
input 	q_b_6;
input 	q_b_7;
input 	q_b_8;
input 	q_b_9;
input 	q_b_10;
input 	q_b_11;
input 	q_b_12;
input 	q_b_13;
input 	q_b_14;
input 	q_b_15;
output 	q_b_01;
output 	q_b_16;
output 	q_b_21;
output 	q_b_31;
output 	q_b_41;
output 	q_b_51;
output 	q_b_61;
output 	q_b_71;
output 	q_b_81;
output 	q_b_91;
output 	q_b_101;
output 	q_b_111;
output 	q_b_121;
output 	q_b_131;
output 	q_b_141;
output 	q_b_151;
input 	always0;
input 	delay_reg_24_0;
input 	short_shift_full;
input 	short_to_long_arrived;
input 	GND_port;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



lms_dsp_altshift_taps_1 ALTSHIFT_TAPS_component(
	.shiftin({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.shiftout({q_b_151,q_b_141,q_b_131,q_b_121,q_b_111,q_b_101,q_b_91,q_b_81,q_b_71,q_b_61,q_b_51,q_b_41,q_b_31,q_b_21,q_b_16,q_b_01}),
	.always0(always0),
	.delay_reg_24_0(delay_reg_24_0),
	.short_shift_full(short_shift_full),
	.clken(short_to_long_arrived),
	.GND_port(GND_port),
	.clock(clk_clk));

endmodule

module lms_dsp_altshift_taps_1 (
	shiftin,
	shiftout,
	always0,
	delay_reg_24_0,
	short_shift_full,
	clken,
	GND_port,
	clock)/* synthesis synthesis_greybox=0 */;
input 	[15:0] shiftin;
output 	[15:0] shiftout;
input 	always0;
input 	delay_reg_24_0;
input 	short_shift_full;
input 	clken;
input 	GND_port;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



lms_dsp_shift_taps_60v auto_generated(
	.shiftin({shiftin[15],shiftin[14],shiftin[13],shiftin[12],shiftin[11],shiftin[10],shiftin[9],shiftin[8],shiftin[7],shiftin[6],shiftin[5],shiftin[4],shiftin[3],shiftin[2],shiftin[1],shiftin[0]}),
	.shiftout({shiftout[15],shiftout[14],shiftout[13],shiftout[12],shiftout[11],shiftout[10],shiftout[9],shiftout[8],shiftout[7],shiftout[6],shiftout[5],shiftout[4],shiftout[3],shiftout[2],shiftout[1],shiftout[0]}),
	.always0(always0),
	.delay_reg_24_0(delay_reg_24_0),
	.short_shift_full(short_shift_full),
	.clken(clken),
	.GND_port(GND_port),
	.clock(clock));

endmodule

module lms_dsp_shift_taps_60v (
	shiftin,
	shiftout,
	always0,
	delay_reg_24_0,
	short_shift_full,
	clken,
	GND_port,
	clock)/* synthesis synthesis_greybox=0 */;
input 	[15:0] shiftin;
output 	[15:0] shiftout;
input 	always0;
input 	delay_reg_24_0;
input 	short_shift_full;
input 	clken;
input 	GND_port;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \cntr1|counter_reg_bit[0]~q ;
wire \cntr1|counter_reg_bit[1]~q ;
wire \cntr1|counter_reg_bit[2]~q ;
wire \cntr1|counter_reg_bit[3]~q ;
wire \cntr1|counter_reg_bit[4]~q ;
wire \cntr1|counter_reg_bit[5]~q ;
wire \cntr1|counter_reg_bit[6]~q ;
wire \cntr1|counter_reg_bit[7]~q ;
wire \cntr3|counter_comb_bita7~0_combout ;
wire \dffe4~q ;


lms_dsp_cntr_0ng cntr3(
	.counter_comb_bita71(\cntr3|counter_comb_bita7~0_combout ),
	.always0(always0),
	.delay_reg_24_0(delay_reg_24_0),
	.short_shift_full(short_shift_full),
	.clock(clock));

lms_dsp_cntr_a7f cntr1(
	.counter_reg_bit_0(\cntr1|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\cntr1|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\cntr1|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\cntr1|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\cntr1|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\cntr1|counter_reg_bit[5]~q ),
	.counter_reg_bit_6(\cntr1|counter_reg_bit[6]~q ),
	.counter_reg_bit_7(\cntr1|counter_reg_bit[7]~q ),
	.short_to_long_arrived(clken),
	.GND_port(GND_port),
	.clock(clock));

lms_dsp_altsyncram_ffc1 altsyncram2(
	.data_a({shiftin[15],shiftin[14],shiftin[13],shiftin[12],shiftin[11],shiftin[10],shiftin[9],shiftin[8],shiftin[7],shiftin[6],shiftin[5],shiftin[4],shiftin[3],shiftin[2],shiftin[1],shiftin[0]}),
	.q_b({shiftout[15],shiftout[14],shiftout[13],shiftout[12],shiftout[11],shiftout[10],shiftout[9],shiftout[8],shiftout[7],shiftout[6],shiftout[5],shiftout[4],shiftout[3],shiftout[2],shiftout[1],shiftout[0]}),
	.address_b({\cntr1|counter_reg_bit[7]~q ,\cntr1|counter_reg_bit[6]~q ,\cntr1|counter_reg_bit[5]~q ,\cntr1|counter_reg_bit[4]~q ,\cntr1|counter_reg_bit[3]~q ,\cntr1|counter_reg_bit[2]~q ,\cntr1|counter_reg_bit[1]~q ,\cntr1|counter_reg_bit[0]~q }),
	.address_a({\cntr1|counter_reg_bit[7]~q ,\cntr1|counter_reg_bit[6]~q ,\cntr1|counter_reg_bit[5]~q ,\cntr1|counter_reg_bit[4]~q ,\cntr1|counter_reg_bit[3]~q ,\cntr1|counter_reg_bit[2]~q ,\cntr1|counter_reg_bit[1]~q ,\cntr1|counter_reg_bit[0]~q }),
	.clocken0(clken),
	.aclr0(\dffe4~q ),
	.clock0(clock));

dffeas dffe4(
	.clk(clock),
	.d(\cntr3|counter_comb_bita7~0_combout ),
	.asdata(vcc),
	.clrn(!always0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dffe4~q ),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

endmodule

module lms_dsp_altsyncram_ffc1 (
	data_a,
	q_b,
	address_b,
	address_a,
	clocken0,
	aclr0,
	clock0)/* synthesis synthesis_greybox=0 */;
input 	[15:0] data_a;
output 	[15:0] q_b;
input 	[7:0] address_b;
input 	[7:0] address_a;
input 	clocken0;
input 	aclr0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block5a0_PORTBDATAOUT_bus;
wire [143:0] ram_block5a1_PORTBDATAOUT_bus;
wire [143:0] ram_block5a2_PORTBDATAOUT_bus;
wire [143:0] ram_block5a3_PORTBDATAOUT_bus;
wire [143:0] ram_block5a4_PORTBDATAOUT_bus;
wire [143:0] ram_block5a5_PORTBDATAOUT_bus;
wire [143:0] ram_block5a6_PORTBDATAOUT_bus;
wire [143:0] ram_block5a7_PORTBDATAOUT_bus;
wire [143:0] ram_block5a8_PORTBDATAOUT_bus;
wire [143:0] ram_block5a9_PORTBDATAOUT_bus;
wire [143:0] ram_block5a10_PORTBDATAOUT_bus;
wire [143:0] ram_block5a11_PORTBDATAOUT_bus;
wire [143:0] ram_block5a12_PORTBDATAOUT_bus;
wire [143:0] ram_block5a13_PORTBDATAOUT_bus;
wire [143:0] ram_block5a14_PORTBDATAOUT_bus;
wire [143:0] ram_block5a15_PORTBDATAOUT_bus;

assign q_b[0] = ram_block5a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block5a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block5a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block5a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block5a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block5a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block5a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block5a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block5a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block5a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block5a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block5a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block5a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block5a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block5a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block5a15_PORTBDATAOUT_bus[0];

fiftyfivenm_ram_block ram_block5a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a0_PORTBDATAOUT_bus));
defparam ram_block5a0.clk0_core_clock_enable = "ena0";
defparam ram_block5a0.clk0_input_clock_enable = "ena0";
defparam ram_block5a0.clk0_output_clock_enable = "ena0";
defparam ram_block5a0.data_interleave_offset_in_bits = 1;
defparam ram_block5a0.data_interleave_width_in_bits = 1;
defparam ram_block5a0.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|long_shift:long_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_60v:auto_generated|altsyncram_ffc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a0.mixed_port_feed_through_mode = "old";
defparam ram_block5a0.operation_mode = "dual_port";
defparam ram_block5a0.port_a_address_clear = "none";
defparam ram_block5a0.port_a_address_width = 8;
defparam ram_block5a0.port_a_data_out_clear = "none";
defparam ram_block5a0.port_a_data_out_clock = "none";
defparam ram_block5a0.port_a_data_width = 1;
defparam ram_block5a0.port_a_first_address = 0;
defparam ram_block5a0.port_a_first_bit_number = 0;
defparam ram_block5a0.port_a_last_address = 253;
defparam ram_block5a0.port_a_logical_ram_depth = 254;
defparam ram_block5a0.port_a_logical_ram_width = 16;
defparam ram_block5a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a0.port_b_address_clear = "none";
defparam ram_block5a0.port_b_address_clock = "clock0";
defparam ram_block5a0.port_b_address_width = 8;
defparam ram_block5a0.port_b_data_out_clear = "clear0";
defparam ram_block5a0.port_b_data_out_clock = "clock0";
defparam ram_block5a0.port_b_data_width = 1;
defparam ram_block5a0.port_b_first_address = 0;
defparam ram_block5a0.port_b_first_bit_number = 0;
defparam ram_block5a0.port_b_last_address = 253;
defparam ram_block5a0.port_b_logical_ram_depth = 254;
defparam ram_block5a0.port_b_logical_ram_width = 16;
defparam ram_block5a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a0.port_b_read_enable_clock = "clock0";
defparam ram_block5a0.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a1_PORTBDATAOUT_bus));
defparam ram_block5a1.clk0_core_clock_enable = "ena0";
defparam ram_block5a1.clk0_input_clock_enable = "ena0";
defparam ram_block5a1.clk0_output_clock_enable = "ena0";
defparam ram_block5a1.data_interleave_offset_in_bits = 1;
defparam ram_block5a1.data_interleave_width_in_bits = 1;
defparam ram_block5a1.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|long_shift:long_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_60v:auto_generated|altsyncram_ffc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a1.mixed_port_feed_through_mode = "old";
defparam ram_block5a1.operation_mode = "dual_port";
defparam ram_block5a1.port_a_address_clear = "none";
defparam ram_block5a1.port_a_address_width = 8;
defparam ram_block5a1.port_a_data_out_clear = "none";
defparam ram_block5a1.port_a_data_out_clock = "none";
defparam ram_block5a1.port_a_data_width = 1;
defparam ram_block5a1.port_a_first_address = 0;
defparam ram_block5a1.port_a_first_bit_number = 1;
defparam ram_block5a1.port_a_last_address = 253;
defparam ram_block5a1.port_a_logical_ram_depth = 254;
defparam ram_block5a1.port_a_logical_ram_width = 16;
defparam ram_block5a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a1.port_b_address_clear = "none";
defparam ram_block5a1.port_b_address_clock = "clock0";
defparam ram_block5a1.port_b_address_width = 8;
defparam ram_block5a1.port_b_data_out_clear = "clear0";
defparam ram_block5a1.port_b_data_out_clock = "clock0";
defparam ram_block5a1.port_b_data_width = 1;
defparam ram_block5a1.port_b_first_address = 0;
defparam ram_block5a1.port_b_first_bit_number = 1;
defparam ram_block5a1.port_b_last_address = 253;
defparam ram_block5a1.port_b_logical_ram_depth = 254;
defparam ram_block5a1.port_b_logical_ram_width = 16;
defparam ram_block5a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a1.port_b_read_enable_clock = "clock0";
defparam ram_block5a1.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a2_PORTBDATAOUT_bus));
defparam ram_block5a2.clk0_core_clock_enable = "ena0";
defparam ram_block5a2.clk0_input_clock_enable = "ena0";
defparam ram_block5a2.clk0_output_clock_enable = "ena0";
defparam ram_block5a2.data_interleave_offset_in_bits = 1;
defparam ram_block5a2.data_interleave_width_in_bits = 1;
defparam ram_block5a2.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|long_shift:long_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_60v:auto_generated|altsyncram_ffc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a2.mixed_port_feed_through_mode = "old";
defparam ram_block5a2.operation_mode = "dual_port";
defparam ram_block5a2.port_a_address_clear = "none";
defparam ram_block5a2.port_a_address_width = 8;
defparam ram_block5a2.port_a_data_out_clear = "none";
defparam ram_block5a2.port_a_data_out_clock = "none";
defparam ram_block5a2.port_a_data_width = 1;
defparam ram_block5a2.port_a_first_address = 0;
defparam ram_block5a2.port_a_first_bit_number = 2;
defparam ram_block5a2.port_a_last_address = 253;
defparam ram_block5a2.port_a_logical_ram_depth = 254;
defparam ram_block5a2.port_a_logical_ram_width = 16;
defparam ram_block5a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a2.port_b_address_clear = "none";
defparam ram_block5a2.port_b_address_clock = "clock0";
defparam ram_block5a2.port_b_address_width = 8;
defparam ram_block5a2.port_b_data_out_clear = "clear0";
defparam ram_block5a2.port_b_data_out_clock = "clock0";
defparam ram_block5a2.port_b_data_width = 1;
defparam ram_block5a2.port_b_first_address = 0;
defparam ram_block5a2.port_b_first_bit_number = 2;
defparam ram_block5a2.port_b_last_address = 253;
defparam ram_block5a2.port_b_logical_ram_depth = 254;
defparam ram_block5a2.port_b_logical_ram_width = 16;
defparam ram_block5a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a2.port_b_read_enable_clock = "clock0";
defparam ram_block5a2.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a3_PORTBDATAOUT_bus));
defparam ram_block5a3.clk0_core_clock_enable = "ena0";
defparam ram_block5a3.clk0_input_clock_enable = "ena0";
defparam ram_block5a3.clk0_output_clock_enable = "ena0";
defparam ram_block5a3.data_interleave_offset_in_bits = 1;
defparam ram_block5a3.data_interleave_width_in_bits = 1;
defparam ram_block5a3.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|long_shift:long_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_60v:auto_generated|altsyncram_ffc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a3.mixed_port_feed_through_mode = "old";
defparam ram_block5a3.operation_mode = "dual_port";
defparam ram_block5a3.port_a_address_clear = "none";
defparam ram_block5a3.port_a_address_width = 8;
defparam ram_block5a3.port_a_data_out_clear = "none";
defparam ram_block5a3.port_a_data_out_clock = "none";
defparam ram_block5a3.port_a_data_width = 1;
defparam ram_block5a3.port_a_first_address = 0;
defparam ram_block5a3.port_a_first_bit_number = 3;
defparam ram_block5a3.port_a_last_address = 253;
defparam ram_block5a3.port_a_logical_ram_depth = 254;
defparam ram_block5a3.port_a_logical_ram_width = 16;
defparam ram_block5a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a3.port_b_address_clear = "none";
defparam ram_block5a3.port_b_address_clock = "clock0";
defparam ram_block5a3.port_b_address_width = 8;
defparam ram_block5a3.port_b_data_out_clear = "clear0";
defparam ram_block5a3.port_b_data_out_clock = "clock0";
defparam ram_block5a3.port_b_data_width = 1;
defparam ram_block5a3.port_b_first_address = 0;
defparam ram_block5a3.port_b_first_bit_number = 3;
defparam ram_block5a3.port_b_last_address = 253;
defparam ram_block5a3.port_b_logical_ram_depth = 254;
defparam ram_block5a3.port_b_logical_ram_width = 16;
defparam ram_block5a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a3.port_b_read_enable_clock = "clock0";
defparam ram_block5a3.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a4_PORTBDATAOUT_bus));
defparam ram_block5a4.clk0_core_clock_enable = "ena0";
defparam ram_block5a4.clk0_input_clock_enable = "ena0";
defparam ram_block5a4.clk0_output_clock_enable = "ena0";
defparam ram_block5a4.data_interleave_offset_in_bits = 1;
defparam ram_block5a4.data_interleave_width_in_bits = 1;
defparam ram_block5a4.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|long_shift:long_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_60v:auto_generated|altsyncram_ffc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a4.mixed_port_feed_through_mode = "old";
defparam ram_block5a4.operation_mode = "dual_port";
defparam ram_block5a4.port_a_address_clear = "none";
defparam ram_block5a4.port_a_address_width = 8;
defparam ram_block5a4.port_a_data_out_clear = "none";
defparam ram_block5a4.port_a_data_out_clock = "none";
defparam ram_block5a4.port_a_data_width = 1;
defparam ram_block5a4.port_a_first_address = 0;
defparam ram_block5a4.port_a_first_bit_number = 4;
defparam ram_block5a4.port_a_last_address = 253;
defparam ram_block5a4.port_a_logical_ram_depth = 254;
defparam ram_block5a4.port_a_logical_ram_width = 16;
defparam ram_block5a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a4.port_b_address_clear = "none";
defparam ram_block5a4.port_b_address_clock = "clock0";
defparam ram_block5a4.port_b_address_width = 8;
defparam ram_block5a4.port_b_data_out_clear = "clear0";
defparam ram_block5a4.port_b_data_out_clock = "clock0";
defparam ram_block5a4.port_b_data_width = 1;
defparam ram_block5a4.port_b_first_address = 0;
defparam ram_block5a4.port_b_first_bit_number = 4;
defparam ram_block5a4.port_b_last_address = 253;
defparam ram_block5a4.port_b_logical_ram_depth = 254;
defparam ram_block5a4.port_b_logical_ram_width = 16;
defparam ram_block5a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a4.port_b_read_enable_clock = "clock0";
defparam ram_block5a4.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a5_PORTBDATAOUT_bus));
defparam ram_block5a5.clk0_core_clock_enable = "ena0";
defparam ram_block5a5.clk0_input_clock_enable = "ena0";
defparam ram_block5a5.clk0_output_clock_enable = "ena0";
defparam ram_block5a5.data_interleave_offset_in_bits = 1;
defparam ram_block5a5.data_interleave_width_in_bits = 1;
defparam ram_block5a5.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|long_shift:long_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_60v:auto_generated|altsyncram_ffc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a5.mixed_port_feed_through_mode = "old";
defparam ram_block5a5.operation_mode = "dual_port";
defparam ram_block5a5.port_a_address_clear = "none";
defparam ram_block5a5.port_a_address_width = 8;
defparam ram_block5a5.port_a_data_out_clear = "none";
defparam ram_block5a5.port_a_data_out_clock = "none";
defparam ram_block5a5.port_a_data_width = 1;
defparam ram_block5a5.port_a_first_address = 0;
defparam ram_block5a5.port_a_first_bit_number = 5;
defparam ram_block5a5.port_a_last_address = 253;
defparam ram_block5a5.port_a_logical_ram_depth = 254;
defparam ram_block5a5.port_a_logical_ram_width = 16;
defparam ram_block5a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a5.port_b_address_clear = "none";
defparam ram_block5a5.port_b_address_clock = "clock0";
defparam ram_block5a5.port_b_address_width = 8;
defparam ram_block5a5.port_b_data_out_clear = "clear0";
defparam ram_block5a5.port_b_data_out_clock = "clock0";
defparam ram_block5a5.port_b_data_width = 1;
defparam ram_block5a5.port_b_first_address = 0;
defparam ram_block5a5.port_b_first_bit_number = 5;
defparam ram_block5a5.port_b_last_address = 253;
defparam ram_block5a5.port_b_logical_ram_depth = 254;
defparam ram_block5a5.port_b_logical_ram_width = 16;
defparam ram_block5a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a5.port_b_read_enable_clock = "clock0";
defparam ram_block5a5.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a6_PORTBDATAOUT_bus));
defparam ram_block5a6.clk0_core_clock_enable = "ena0";
defparam ram_block5a6.clk0_input_clock_enable = "ena0";
defparam ram_block5a6.clk0_output_clock_enable = "ena0";
defparam ram_block5a6.data_interleave_offset_in_bits = 1;
defparam ram_block5a6.data_interleave_width_in_bits = 1;
defparam ram_block5a6.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|long_shift:long_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_60v:auto_generated|altsyncram_ffc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a6.mixed_port_feed_through_mode = "old";
defparam ram_block5a6.operation_mode = "dual_port";
defparam ram_block5a6.port_a_address_clear = "none";
defparam ram_block5a6.port_a_address_width = 8;
defparam ram_block5a6.port_a_data_out_clear = "none";
defparam ram_block5a6.port_a_data_out_clock = "none";
defparam ram_block5a6.port_a_data_width = 1;
defparam ram_block5a6.port_a_first_address = 0;
defparam ram_block5a6.port_a_first_bit_number = 6;
defparam ram_block5a6.port_a_last_address = 253;
defparam ram_block5a6.port_a_logical_ram_depth = 254;
defparam ram_block5a6.port_a_logical_ram_width = 16;
defparam ram_block5a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a6.port_b_address_clear = "none";
defparam ram_block5a6.port_b_address_clock = "clock0";
defparam ram_block5a6.port_b_address_width = 8;
defparam ram_block5a6.port_b_data_out_clear = "clear0";
defparam ram_block5a6.port_b_data_out_clock = "clock0";
defparam ram_block5a6.port_b_data_width = 1;
defparam ram_block5a6.port_b_first_address = 0;
defparam ram_block5a6.port_b_first_bit_number = 6;
defparam ram_block5a6.port_b_last_address = 253;
defparam ram_block5a6.port_b_logical_ram_depth = 254;
defparam ram_block5a6.port_b_logical_ram_width = 16;
defparam ram_block5a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a6.port_b_read_enable_clock = "clock0";
defparam ram_block5a6.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a7_PORTBDATAOUT_bus));
defparam ram_block5a7.clk0_core_clock_enable = "ena0";
defparam ram_block5a7.clk0_input_clock_enable = "ena0";
defparam ram_block5a7.clk0_output_clock_enable = "ena0";
defparam ram_block5a7.data_interleave_offset_in_bits = 1;
defparam ram_block5a7.data_interleave_width_in_bits = 1;
defparam ram_block5a7.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|long_shift:long_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_60v:auto_generated|altsyncram_ffc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a7.mixed_port_feed_through_mode = "old";
defparam ram_block5a7.operation_mode = "dual_port";
defparam ram_block5a7.port_a_address_clear = "none";
defparam ram_block5a7.port_a_address_width = 8;
defparam ram_block5a7.port_a_data_out_clear = "none";
defparam ram_block5a7.port_a_data_out_clock = "none";
defparam ram_block5a7.port_a_data_width = 1;
defparam ram_block5a7.port_a_first_address = 0;
defparam ram_block5a7.port_a_first_bit_number = 7;
defparam ram_block5a7.port_a_last_address = 253;
defparam ram_block5a7.port_a_logical_ram_depth = 254;
defparam ram_block5a7.port_a_logical_ram_width = 16;
defparam ram_block5a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a7.port_b_address_clear = "none";
defparam ram_block5a7.port_b_address_clock = "clock0";
defparam ram_block5a7.port_b_address_width = 8;
defparam ram_block5a7.port_b_data_out_clear = "clear0";
defparam ram_block5a7.port_b_data_out_clock = "clock0";
defparam ram_block5a7.port_b_data_width = 1;
defparam ram_block5a7.port_b_first_address = 0;
defparam ram_block5a7.port_b_first_bit_number = 7;
defparam ram_block5a7.port_b_last_address = 253;
defparam ram_block5a7.port_b_logical_ram_depth = 254;
defparam ram_block5a7.port_b_logical_ram_width = 16;
defparam ram_block5a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a7.port_b_read_enable_clock = "clock0";
defparam ram_block5a7.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a8(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a8_PORTBDATAOUT_bus));
defparam ram_block5a8.clk0_core_clock_enable = "ena0";
defparam ram_block5a8.clk0_input_clock_enable = "ena0";
defparam ram_block5a8.clk0_output_clock_enable = "ena0";
defparam ram_block5a8.data_interleave_offset_in_bits = 1;
defparam ram_block5a8.data_interleave_width_in_bits = 1;
defparam ram_block5a8.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|long_shift:long_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_60v:auto_generated|altsyncram_ffc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a8.mixed_port_feed_through_mode = "old";
defparam ram_block5a8.operation_mode = "dual_port";
defparam ram_block5a8.port_a_address_clear = "none";
defparam ram_block5a8.port_a_address_width = 8;
defparam ram_block5a8.port_a_data_out_clear = "none";
defparam ram_block5a8.port_a_data_out_clock = "none";
defparam ram_block5a8.port_a_data_width = 1;
defparam ram_block5a8.port_a_first_address = 0;
defparam ram_block5a8.port_a_first_bit_number = 8;
defparam ram_block5a8.port_a_last_address = 253;
defparam ram_block5a8.port_a_logical_ram_depth = 254;
defparam ram_block5a8.port_a_logical_ram_width = 16;
defparam ram_block5a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a8.port_b_address_clear = "none";
defparam ram_block5a8.port_b_address_clock = "clock0";
defparam ram_block5a8.port_b_address_width = 8;
defparam ram_block5a8.port_b_data_out_clear = "clear0";
defparam ram_block5a8.port_b_data_out_clock = "clock0";
defparam ram_block5a8.port_b_data_width = 1;
defparam ram_block5a8.port_b_first_address = 0;
defparam ram_block5a8.port_b_first_bit_number = 8;
defparam ram_block5a8.port_b_last_address = 253;
defparam ram_block5a8.port_b_logical_ram_depth = 254;
defparam ram_block5a8.port_b_logical_ram_width = 16;
defparam ram_block5a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a8.port_b_read_enable_clock = "clock0";
defparam ram_block5a8.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a9(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a9_PORTBDATAOUT_bus));
defparam ram_block5a9.clk0_core_clock_enable = "ena0";
defparam ram_block5a9.clk0_input_clock_enable = "ena0";
defparam ram_block5a9.clk0_output_clock_enable = "ena0";
defparam ram_block5a9.data_interleave_offset_in_bits = 1;
defparam ram_block5a9.data_interleave_width_in_bits = 1;
defparam ram_block5a9.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|long_shift:long_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_60v:auto_generated|altsyncram_ffc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a9.mixed_port_feed_through_mode = "old";
defparam ram_block5a9.operation_mode = "dual_port";
defparam ram_block5a9.port_a_address_clear = "none";
defparam ram_block5a9.port_a_address_width = 8;
defparam ram_block5a9.port_a_data_out_clear = "none";
defparam ram_block5a9.port_a_data_out_clock = "none";
defparam ram_block5a9.port_a_data_width = 1;
defparam ram_block5a9.port_a_first_address = 0;
defparam ram_block5a9.port_a_first_bit_number = 9;
defparam ram_block5a9.port_a_last_address = 253;
defparam ram_block5a9.port_a_logical_ram_depth = 254;
defparam ram_block5a9.port_a_logical_ram_width = 16;
defparam ram_block5a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a9.port_b_address_clear = "none";
defparam ram_block5a9.port_b_address_clock = "clock0";
defparam ram_block5a9.port_b_address_width = 8;
defparam ram_block5a9.port_b_data_out_clear = "clear0";
defparam ram_block5a9.port_b_data_out_clock = "clock0";
defparam ram_block5a9.port_b_data_width = 1;
defparam ram_block5a9.port_b_first_address = 0;
defparam ram_block5a9.port_b_first_bit_number = 9;
defparam ram_block5a9.port_b_last_address = 253;
defparam ram_block5a9.port_b_logical_ram_depth = 254;
defparam ram_block5a9.port_b_logical_ram_width = 16;
defparam ram_block5a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a9.port_b_read_enable_clock = "clock0";
defparam ram_block5a9.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a10(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a10_PORTBDATAOUT_bus));
defparam ram_block5a10.clk0_core_clock_enable = "ena0";
defparam ram_block5a10.clk0_input_clock_enable = "ena0";
defparam ram_block5a10.clk0_output_clock_enable = "ena0";
defparam ram_block5a10.data_interleave_offset_in_bits = 1;
defparam ram_block5a10.data_interleave_width_in_bits = 1;
defparam ram_block5a10.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|long_shift:long_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_60v:auto_generated|altsyncram_ffc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a10.mixed_port_feed_through_mode = "old";
defparam ram_block5a10.operation_mode = "dual_port";
defparam ram_block5a10.port_a_address_clear = "none";
defparam ram_block5a10.port_a_address_width = 8;
defparam ram_block5a10.port_a_data_out_clear = "none";
defparam ram_block5a10.port_a_data_out_clock = "none";
defparam ram_block5a10.port_a_data_width = 1;
defparam ram_block5a10.port_a_first_address = 0;
defparam ram_block5a10.port_a_first_bit_number = 10;
defparam ram_block5a10.port_a_last_address = 253;
defparam ram_block5a10.port_a_logical_ram_depth = 254;
defparam ram_block5a10.port_a_logical_ram_width = 16;
defparam ram_block5a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a10.port_b_address_clear = "none";
defparam ram_block5a10.port_b_address_clock = "clock0";
defparam ram_block5a10.port_b_address_width = 8;
defparam ram_block5a10.port_b_data_out_clear = "clear0";
defparam ram_block5a10.port_b_data_out_clock = "clock0";
defparam ram_block5a10.port_b_data_width = 1;
defparam ram_block5a10.port_b_first_address = 0;
defparam ram_block5a10.port_b_first_bit_number = 10;
defparam ram_block5a10.port_b_last_address = 253;
defparam ram_block5a10.port_b_logical_ram_depth = 254;
defparam ram_block5a10.port_b_logical_ram_width = 16;
defparam ram_block5a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a10.port_b_read_enable_clock = "clock0";
defparam ram_block5a10.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a11(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a11_PORTBDATAOUT_bus));
defparam ram_block5a11.clk0_core_clock_enable = "ena0";
defparam ram_block5a11.clk0_input_clock_enable = "ena0";
defparam ram_block5a11.clk0_output_clock_enable = "ena0";
defparam ram_block5a11.data_interleave_offset_in_bits = 1;
defparam ram_block5a11.data_interleave_width_in_bits = 1;
defparam ram_block5a11.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|long_shift:long_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_60v:auto_generated|altsyncram_ffc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a11.mixed_port_feed_through_mode = "old";
defparam ram_block5a11.operation_mode = "dual_port";
defparam ram_block5a11.port_a_address_clear = "none";
defparam ram_block5a11.port_a_address_width = 8;
defparam ram_block5a11.port_a_data_out_clear = "none";
defparam ram_block5a11.port_a_data_out_clock = "none";
defparam ram_block5a11.port_a_data_width = 1;
defparam ram_block5a11.port_a_first_address = 0;
defparam ram_block5a11.port_a_first_bit_number = 11;
defparam ram_block5a11.port_a_last_address = 253;
defparam ram_block5a11.port_a_logical_ram_depth = 254;
defparam ram_block5a11.port_a_logical_ram_width = 16;
defparam ram_block5a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a11.port_b_address_clear = "none";
defparam ram_block5a11.port_b_address_clock = "clock0";
defparam ram_block5a11.port_b_address_width = 8;
defparam ram_block5a11.port_b_data_out_clear = "clear0";
defparam ram_block5a11.port_b_data_out_clock = "clock0";
defparam ram_block5a11.port_b_data_width = 1;
defparam ram_block5a11.port_b_first_address = 0;
defparam ram_block5a11.port_b_first_bit_number = 11;
defparam ram_block5a11.port_b_last_address = 253;
defparam ram_block5a11.port_b_logical_ram_depth = 254;
defparam ram_block5a11.port_b_logical_ram_width = 16;
defparam ram_block5a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a11.port_b_read_enable_clock = "clock0";
defparam ram_block5a11.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a12(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a12_PORTBDATAOUT_bus));
defparam ram_block5a12.clk0_core_clock_enable = "ena0";
defparam ram_block5a12.clk0_input_clock_enable = "ena0";
defparam ram_block5a12.clk0_output_clock_enable = "ena0";
defparam ram_block5a12.data_interleave_offset_in_bits = 1;
defparam ram_block5a12.data_interleave_width_in_bits = 1;
defparam ram_block5a12.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|long_shift:long_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_60v:auto_generated|altsyncram_ffc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a12.mixed_port_feed_through_mode = "old";
defparam ram_block5a12.operation_mode = "dual_port";
defparam ram_block5a12.port_a_address_clear = "none";
defparam ram_block5a12.port_a_address_width = 8;
defparam ram_block5a12.port_a_data_out_clear = "none";
defparam ram_block5a12.port_a_data_out_clock = "none";
defparam ram_block5a12.port_a_data_width = 1;
defparam ram_block5a12.port_a_first_address = 0;
defparam ram_block5a12.port_a_first_bit_number = 12;
defparam ram_block5a12.port_a_last_address = 253;
defparam ram_block5a12.port_a_logical_ram_depth = 254;
defparam ram_block5a12.port_a_logical_ram_width = 16;
defparam ram_block5a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a12.port_b_address_clear = "none";
defparam ram_block5a12.port_b_address_clock = "clock0";
defparam ram_block5a12.port_b_address_width = 8;
defparam ram_block5a12.port_b_data_out_clear = "clear0";
defparam ram_block5a12.port_b_data_out_clock = "clock0";
defparam ram_block5a12.port_b_data_width = 1;
defparam ram_block5a12.port_b_first_address = 0;
defparam ram_block5a12.port_b_first_bit_number = 12;
defparam ram_block5a12.port_b_last_address = 253;
defparam ram_block5a12.port_b_logical_ram_depth = 254;
defparam ram_block5a12.port_b_logical_ram_width = 16;
defparam ram_block5a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a12.port_b_read_enable_clock = "clock0";
defparam ram_block5a12.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a13(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a13_PORTBDATAOUT_bus));
defparam ram_block5a13.clk0_core_clock_enable = "ena0";
defparam ram_block5a13.clk0_input_clock_enable = "ena0";
defparam ram_block5a13.clk0_output_clock_enable = "ena0";
defparam ram_block5a13.data_interleave_offset_in_bits = 1;
defparam ram_block5a13.data_interleave_width_in_bits = 1;
defparam ram_block5a13.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|long_shift:long_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_60v:auto_generated|altsyncram_ffc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a13.mixed_port_feed_through_mode = "old";
defparam ram_block5a13.operation_mode = "dual_port";
defparam ram_block5a13.port_a_address_clear = "none";
defparam ram_block5a13.port_a_address_width = 8;
defparam ram_block5a13.port_a_data_out_clear = "none";
defparam ram_block5a13.port_a_data_out_clock = "none";
defparam ram_block5a13.port_a_data_width = 1;
defparam ram_block5a13.port_a_first_address = 0;
defparam ram_block5a13.port_a_first_bit_number = 13;
defparam ram_block5a13.port_a_last_address = 253;
defparam ram_block5a13.port_a_logical_ram_depth = 254;
defparam ram_block5a13.port_a_logical_ram_width = 16;
defparam ram_block5a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a13.port_b_address_clear = "none";
defparam ram_block5a13.port_b_address_clock = "clock0";
defparam ram_block5a13.port_b_address_width = 8;
defparam ram_block5a13.port_b_data_out_clear = "clear0";
defparam ram_block5a13.port_b_data_out_clock = "clock0";
defparam ram_block5a13.port_b_data_width = 1;
defparam ram_block5a13.port_b_first_address = 0;
defparam ram_block5a13.port_b_first_bit_number = 13;
defparam ram_block5a13.port_b_last_address = 253;
defparam ram_block5a13.port_b_logical_ram_depth = 254;
defparam ram_block5a13.port_b_logical_ram_width = 16;
defparam ram_block5a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a13.port_b_read_enable_clock = "clock0";
defparam ram_block5a13.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a14(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a14_PORTBDATAOUT_bus));
defparam ram_block5a14.clk0_core_clock_enable = "ena0";
defparam ram_block5a14.clk0_input_clock_enable = "ena0";
defparam ram_block5a14.clk0_output_clock_enable = "ena0";
defparam ram_block5a14.data_interleave_offset_in_bits = 1;
defparam ram_block5a14.data_interleave_width_in_bits = 1;
defparam ram_block5a14.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|long_shift:long_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_60v:auto_generated|altsyncram_ffc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a14.mixed_port_feed_through_mode = "old";
defparam ram_block5a14.operation_mode = "dual_port";
defparam ram_block5a14.port_a_address_clear = "none";
defparam ram_block5a14.port_a_address_width = 8;
defparam ram_block5a14.port_a_data_out_clear = "none";
defparam ram_block5a14.port_a_data_out_clock = "none";
defparam ram_block5a14.port_a_data_width = 1;
defparam ram_block5a14.port_a_first_address = 0;
defparam ram_block5a14.port_a_first_bit_number = 14;
defparam ram_block5a14.port_a_last_address = 253;
defparam ram_block5a14.port_a_logical_ram_depth = 254;
defparam ram_block5a14.port_a_logical_ram_width = 16;
defparam ram_block5a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a14.port_b_address_clear = "none";
defparam ram_block5a14.port_b_address_clock = "clock0";
defparam ram_block5a14.port_b_address_width = 8;
defparam ram_block5a14.port_b_data_out_clear = "clear0";
defparam ram_block5a14.port_b_data_out_clock = "clock0";
defparam ram_block5a14.port_b_data_width = 1;
defparam ram_block5a14.port_b_first_address = 0;
defparam ram_block5a14.port_b_first_bit_number = 14;
defparam ram_block5a14.port_b_last_address = 253;
defparam ram_block5a14.port_b_logical_ram_depth = 254;
defparam ram_block5a14.port_b_logical_ram_width = 16;
defparam ram_block5a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a14.port_b_read_enable_clock = "clock0";
defparam ram_block5a14.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a15(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a15_PORTBDATAOUT_bus));
defparam ram_block5a15.clk0_core_clock_enable = "ena0";
defparam ram_block5a15.clk0_input_clock_enable = "ena0";
defparam ram_block5a15.clk0_output_clock_enable = "ena0";
defparam ram_block5a15.data_interleave_offset_in_bits = 1;
defparam ram_block5a15.data_interleave_width_in_bits = 1;
defparam ram_block5a15.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|long_shift:long_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_60v:auto_generated|altsyncram_ffc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a15.mixed_port_feed_through_mode = "old";
defparam ram_block5a15.operation_mode = "dual_port";
defparam ram_block5a15.port_a_address_clear = "none";
defparam ram_block5a15.port_a_address_width = 8;
defparam ram_block5a15.port_a_data_out_clear = "none";
defparam ram_block5a15.port_a_data_out_clock = "none";
defparam ram_block5a15.port_a_data_width = 1;
defparam ram_block5a15.port_a_first_address = 0;
defparam ram_block5a15.port_a_first_bit_number = 15;
defparam ram_block5a15.port_a_last_address = 253;
defparam ram_block5a15.port_a_logical_ram_depth = 254;
defparam ram_block5a15.port_a_logical_ram_width = 16;
defparam ram_block5a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a15.port_b_address_clear = "none";
defparam ram_block5a15.port_b_address_clock = "clock0";
defparam ram_block5a15.port_b_address_width = 8;
defparam ram_block5a15.port_b_data_out_clear = "clear0";
defparam ram_block5a15.port_b_data_out_clock = "clock0";
defparam ram_block5a15.port_b_data_width = 1;
defparam ram_block5a15.port_b_first_address = 0;
defparam ram_block5a15.port_b_first_bit_number = 15;
defparam ram_block5a15.port_b_last_address = 253;
defparam ram_block5a15.port_b_logical_ram_depth = 254;
defparam ram_block5a15.port_b_logical_ram_width = 16;
defparam ram_block5a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a15.port_b_read_enable_clock = "clock0";
defparam ram_block5a15.ram_block_type = "M9K";

endmodule

module lms_dsp_cntr_0ng (
	counter_comb_bita71,
	always0,
	delay_reg_24_0,
	short_shift_full,
	clock)/* synthesis synthesis_greybox=0 */;
output 	counter_comb_bita71;
input 	always0;
input 	delay_reg_24_0;
input 	short_shift_full;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_reg_bit[7]~2_combout ;
wire \counter_reg_bit[0]~q ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_reg_bit[1]~q ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_reg_bit[2]~q ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_reg_bit[3]~q ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_reg_bit[4]~q ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_reg_bit[5]~q ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~combout ;
wire \counter_reg_bit[6]~q ;
wire \counter_comb_bita6~COUT ;
wire \counter_comb_bita7~combout ;
wire \counter_reg_bit[7]~q ;
wire \counter_comb_bita7~COUT ;


fiftyfivenm_lcell_comb \counter_comb_bita7~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita7~COUT ),
	.combout(counter_comb_bita71),
	.cout());
defparam \counter_comb_bita7~0 .lut_mask = 16'h0F0F;
defparam \counter_comb_bita7~0 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(\counter_reg_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5555;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter_reg_bit[7]~2 (
	.dataa(delay_reg_24_0),
	.datab(short_shift_full),
	.datac(counter_comb_bita71),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter_reg_bit[7]~2_combout ),
	.cout());
defparam \counter_reg_bit[7]~2 .lut_mask = 16'h0808;
defparam \counter_reg_bit[7]~2 .sum_lutc_input = "datac";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!always0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\counter_reg_bit[7]~2_combout ),
	.q(\counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(\counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!always0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\counter_reg_bit[7]~2_combout ),
	.q(\counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(\counter_reg_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'hA50A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!always0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\counter_reg_bit[7]~2_combout ),
	.q(\counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(\counter_reg_bit[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!always0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\counter_reg_bit[7]~2_combout ),
	.q(\counter_reg_bit[3]~q ),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita4(
	.dataa(\counter_reg_bit[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'hA50A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!always0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\counter_reg_bit[7]~2_combout ),
	.q(\counter_reg_bit[4]~q ),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita5(
	.dataa(\counter_reg_bit[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout(\counter_comb_bita5~COUT ));
defparam counter_comb_bita5.lut_mask = 16'h5A5F;
defparam counter_comb_bita5.sum_lutc_input = "cin";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!always0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\counter_reg_bit[7]~2_combout ),
	.q(\counter_reg_bit[5]~q ),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita6(
	.dataa(\counter_reg_bit[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita5~COUT ),
	.combout(\counter_comb_bita6~combout ),
	.cout(\counter_comb_bita6~COUT ));
defparam counter_comb_bita6.lut_mask = 16'hA50A;
defparam counter_comb_bita6.sum_lutc_input = "cin";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~combout ),
	.asdata(vcc),
	.clrn(!always0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\counter_reg_bit[7]~2_combout ),
	.q(\counter_reg_bit[6]~q ),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita7(
	.dataa(\counter_reg_bit[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita6~COUT ),
	.combout(\counter_comb_bita7~combout ),
	.cout(\counter_comb_bita7~COUT ));
defparam counter_comb_bita7.lut_mask = 16'h5A5F;
defparam counter_comb_bita7.sum_lutc_input = "cin";

dffeas \counter_reg_bit[7] (
	.clk(clock),
	.d(\counter_comb_bita7~combout ),
	.asdata(vcc),
	.clrn(!always0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\counter_reg_bit[7]~2_combout ),
	.q(\counter_reg_bit[7]~q ),
	.prn(vcc));
defparam \counter_reg_bit[7] .is_wysiwyg = "true";
defparam \counter_reg_bit[7] .power_up = "low";

endmodule

module lms_dsp_cntr_a7f (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	counter_reg_bit_6,
	counter_reg_bit_7,
	short_to_long_arrived,
	GND_port,
	clock)/* synthesis synthesis_greybox=0 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
output 	counter_reg_bit_6;
output 	counter_reg_bit_7;
input 	short_to_long_arrived;
input 	GND_port;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \cmpr6|aneb_result_wire[0]~0_combout ;
wire \cmpr6|aneb_result_wire[0]~1_combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~COUT ;
wire \counter_comb_bita7~COUT ;
wire \counter_comb_bita7~0_combout ;
wire \cout_actual~combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita6~combout ;
wire \counter_comb_bita7~combout ;


lms_dsp_cmpr_krb cmpr6(
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_7(counter_reg_bit_7),
	.aneb_result_wire_0(\cmpr6|aneb_result_wire[0]~0_combout ),
	.aneb_result_wire_01(\cmpr6|aneb_result_wire[0]~1_combout ));

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\cout_actual~combout ),
	.ena(short_to_long_arrived),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\cout_actual~combout ),
	.ena(short_to_long_arrived),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\cout_actual~combout ),
	.ena(short_to_long_arrived),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\cout_actual~combout ),
	.ena(short_to_long_arrived),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\cout_actual~combout ),
	.ena(short_to_long_arrived),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\cout_actual~combout ),
	.ena(short_to_long_arrived),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\cout_actual~combout ),
	.ena(short_to_long_arrived),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

dffeas \counter_reg_bit[7] (
	.clk(clock),
	.d(\counter_comb_bita7~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\cout_actual~combout ),
	.ena(short_to_long_arrived),
	.q(counter_reg_bit_7),
	.prn(vcc));
defparam \counter_reg_bit[7] .is_wysiwyg = "true";
defparam \counter_reg_bit[7] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'hA50A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'hA50A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout(\counter_comb_bita5~COUT ));
defparam counter_comb_bita5.lut_mask = 16'h5A5F;
defparam counter_comb_bita5.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita6(
	.dataa(counter_reg_bit_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita5~COUT ),
	.combout(\counter_comb_bita6~combout ),
	.cout(\counter_comb_bita6~COUT ));
defparam counter_comb_bita6.lut_mask = 16'hA50A;
defparam counter_comb_bita6.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita7(
	.dataa(counter_reg_bit_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita6~COUT ),
	.combout(\counter_comb_bita7~combout ),
	.cout(\counter_comb_bita7~COUT ));
defparam counter_comb_bita7.lut_mask = 16'h5A5F;
defparam counter_comb_bita7.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter_comb_bita7~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita7~COUT ),
	.combout(\counter_comb_bita7~0_combout ),
	.cout());
defparam \counter_comb_bita7~0 .lut_mask = 16'h0F0F;
defparam \counter_comb_bita7~0 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb cout_actual(
	.dataa(\counter_comb_bita7~0_combout ),
	.datab(\cmpr6|aneb_result_wire[0]~0_combout ),
	.datac(\cmpr6|aneb_result_wire[0]~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\cout_actual~combout ),
	.cout());
defparam cout_actual.lut_mask = 16'hEAEA;
defparam cout_actual.sum_lutc_input = "datac";

endmodule

module lms_dsp_cmpr_krb (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	counter_reg_bit_6,
	counter_reg_bit_7,
	aneb_result_wire_0,
	aneb_result_wire_01)/* synthesis synthesis_greybox=0 */;
input 	counter_reg_bit_0;
input 	counter_reg_bit_1;
input 	counter_reg_bit_2;
input 	counter_reg_bit_3;
input 	counter_reg_bit_4;
input 	counter_reg_bit_5;
input 	counter_reg_bit_6;
input 	counter_reg_bit_7;
output 	aneb_result_wire_0;
output 	aneb_result_wire_01;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fiftyfivenm_lcell_comb \aneb_result_wire[0]~0 (
	.dataa(counter_reg_bit_4),
	.datab(counter_reg_bit_5),
	.datac(counter_reg_bit_6),
	.datad(counter_reg_bit_7),
	.cin(gnd),
	.combout(aneb_result_wire_0),
	.cout());
defparam \aneb_result_wire[0]~0 .lut_mask = 16'h8000;
defparam \aneb_result_wire[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \aneb_result_wire[0]~1 (
	.dataa(counter_reg_bit_0),
	.datab(counter_reg_bit_2),
	.datac(counter_reg_bit_3),
	.datad(counter_reg_bit_1),
	.cin(gnd),
	.combout(aneb_result_wire_01),
	.cout());
defparam \aneb_result_wire[0]~1 .lut_mask = 16'h0080;
defparam \aneb_result_wire[0]~1 .sum_lutc_input = "datac";

endmodule

module lms_dsp_short_shift (
	mag_reg_0,
	q_b_0,
	mag_reg_1,
	q_b_1,
	mag_reg_2,
	q_b_2,
	mag_reg_3,
	q_b_3,
	mag_reg_4,
	q_b_4,
	mag_reg_5,
	q_b_5,
	mag_reg_6,
	q_b_6,
	mag_reg_7,
	q_b_7,
	mag_reg_8,
	q_b_8,
	mag_reg_9,
	q_b_9,
	mag_reg_10,
	q_b_10,
	mag_reg_11,
	q_b_11,
	mag_reg_12,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	always0,
	delay_reg_24_0,
	GND_port,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	mag_reg_0;
output 	q_b_0;
input 	mag_reg_1;
output 	q_b_1;
input 	mag_reg_2;
output 	q_b_2;
input 	mag_reg_3;
output 	q_b_3;
input 	mag_reg_4;
output 	q_b_4;
input 	mag_reg_5;
output 	q_b_5;
input 	mag_reg_6;
output 	q_b_6;
input 	mag_reg_7;
output 	q_b_7;
input 	mag_reg_8;
output 	q_b_8;
input 	mag_reg_9;
output 	q_b_9;
input 	mag_reg_10;
output 	q_b_10;
input 	mag_reg_11;
output 	q_b_11;
input 	mag_reg_12;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
input 	always0;
input 	delay_reg_24_0;
input 	GND_port;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



lms_dsp_altshift_taps_2 ALTSHIFT_TAPS_component(
	.shiftin({gnd,gnd,GND_port,mag_reg_12,mag_reg_11,mag_reg_10,mag_reg_9,mag_reg_8,mag_reg_7,mag_reg_6,mag_reg_5,mag_reg_4,mag_reg_3,mag_reg_2,mag_reg_1,mag_reg_0}),
	.shiftout({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.always0(always0),
	.clken(delay_reg_24_0),
	.clock(clk_clk));

endmodule

module lms_dsp_altshift_taps_2 (
	shiftin,
	shiftout,
	always0,
	clken,
	clock)/* synthesis synthesis_greybox=0 */;
input 	[15:0] shiftin;
output 	[15:0] shiftout;
input 	always0;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



lms_dsp_shift_taps_euu auto_generated(
	.shiftin({gnd,gnd,shiftin[13],shiftin[12],shiftin[11],shiftin[10],shiftin[9],shiftin[8],shiftin[7],shiftin[6],shiftin[5],shiftin[4],shiftin[3],shiftin[2],shiftin[1],shiftin[0]}),
	.shiftout({shiftout[15],shiftout[14],shiftout[13],shiftout[12],shiftout[11],shiftout[10],shiftout[9],shiftout[8],shiftout[7],shiftout[6],shiftout[5],shiftout[4],shiftout[3],shiftout[2],shiftout[1],shiftout[0]}),
	.always0(always0),
	.clken(clken),
	.clock(clock));

endmodule

module lms_dsp_shift_taps_euu (
	shiftin,
	shiftout,
	always0,
	clken,
	clock)/* synthesis synthesis_greybox=0 */;
input 	[15:0] shiftin;
output 	[15:0] shiftout;
input 	always0;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \cntr1|counter_reg_bit[0]~q ;
wire \cntr1|counter_reg_bit[1]~q ;
wire \cntr1|counter_reg_bit[2]~q ;
wire \cntr1|counter_reg_bit[3]~q ;
wire \cntr1|counter_reg_bit[4]~q ;
wire \cntr3|counter_comb_bita4~0_combout ;
wire \dffe4~q ;


lms_dsp_cntr_5lg cntr3(
	.counter_comb_bita41(\cntr3|counter_comb_bita4~0_combout ),
	.always0(always0),
	.delay_reg_24_0(clken),
	.clock(clock));

lms_dsp_cntr_f5f cntr1(
	.counter_reg_bit_0(\cntr1|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\cntr1|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\cntr1|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\cntr1|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\cntr1|counter_reg_bit[4]~q ),
	.delay_reg_24_0(clken),
	.GND_port(shiftin[13]),
	.clock(clock));

lms_dsp_altsyncram_pbc1 altsyncram2(
	.data_a({shiftin[13],shiftin[13],shiftin[13],shiftin[12],shiftin[11],shiftin[10],shiftin[9],shiftin[8],shiftin[7],shiftin[6],shiftin[5],shiftin[4],shiftin[3],shiftin[2],shiftin[1],shiftin[0]}),
	.q_b({shiftout[15],shiftout[14],shiftout[13],shiftout[12],shiftout[11],shiftout[10],shiftout[9],shiftout[8],shiftout[7],shiftout[6],shiftout[5],shiftout[4],shiftout[3],shiftout[2],shiftout[1],shiftout[0]}),
	.address_b({\cntr1|counter_reg_bit[4]~q ,\cntr1|counter_reg_bit[3]~q ,\cntr1|counter_reg_bit[2]~q ,\cntr1|counter_reg_bit[1]~q ,\cntr1|counter_reg_bit[0]~q }),
	.address_a({\cntr1|counter_reg_bit[4]~q ,\cntr1|counter_reg_bit[3]~q ,\cntr1|counter_reg_bit[2]~q ,\cntr1|counter_reg_bit[1]~q ,\cntr1|counter_reg_bit[0]~q }),
	.clocken0(clken),
	.aclr0(\dffe4~q ),
	.clock0(clock));

dffeas dffe4(
	.clk(clock),
	.d(\cntr3|counter_comb_bita4~0_combout ),
	.asdata(vcc),
	.clrn(!always0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dffe4~q ),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

endmodule

module lms_dsp_altsyncram_pbc1 (
	data_a,
	q_b,
	address_b,
	address_a,
	clocken0,
	aclr0,
	clock0)/* synthesis synthesis_greybox=0 */;
input 	[15:0] data_a;
output 	[15:0] q_b;
input 	[4:0] address_b;
input 	[4:0] address_a;
input 	clocken0;
input 	aclr0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block5a0_PORTBDATAOUT_bus;
wire [143:0] ram_block5a1_PORTBDATAOUT_bus;
wire [143:0] ram_block5a2_PORTBDATAOUT_bus;
wire [143:0] ram_block5a3_PORTBDATAOUT_bus;
wire [143:0] ram_block5a4_PORTBDATAOUT_bus;
wire [143:0] ram_block5a5_PORTBDATAOUT_bus;
wire [143:0] ram_block5a6_PORTBDATAOUT_bus;
wire [143:0] ram_block5a7_PORTBDATAOUT_bus;
wire [143:0] ram_block5a8_PORTBDATAOUT_bus;
wire [143:0] ram_block5a9_PORTBDATAOUT_bus;
wire [143:0] ram_block5a10_PORTBDATAOUT_bus;
wire [143:0] ram_block5a11_PORTBDATAOUT_bus;
wire [143:0] ram_block5a12_PORTBDATAOUT_bus;
wire [143:0] ram_block5a13_PORTBDATAOUT_bus;
wire [143:0] ram_block5a14_PORTBDATAOUT_bus;
wire [143:0] ram_block5a15_PORTBDATAOUT_bus;

assign q_b[0] = ram_block5a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block5a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block5a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block5a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block5a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block5a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block5a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block5a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block5a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block5a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block5a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block5a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block5a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block5a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block5a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block5a15_PORTBDATAOUT_bus[0];

fiftyfivenm_ram_block ram_block5a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a0_PORTBDATAOUT_bus));
defparam ram_block5a0.clk0_core_clock_enable = "ena0";
defparam ram_block5a0.clk0_input_clock_enable = "ena0";
defparam ram_block5a0.clk0_output_clock_enable = "ena0";
defparam ram_block5a0.data_interleave_offset_in_bits = 1;
defparam ram_block5a0.data_interleave_width_in_bits = 1;
defparam ram_block5a0.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|short_shift:short_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_euu:auto_generated|altsyncram_pbc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a0.mixed_port_feed_through_mode = "old";
defparam ram_block5a0.operation_mode = "dual_port";
defparam ram_block5a0.port_a_address_clear = "none";
defparam ram_block5a0.port_a_address_width = 5;
defparam ram_block5a0.port_a_data_out_clear = "none";
defparam ram_block5a0.port_a_data_out_clock = "none";
defparam ram_block5a0.port_a_data_width = 1;
defparam ram_block5a0.port_a_first_address = 0;
defparam ram_block5a0.port_a_first_bit_number = 0;
defparam ram_block5a0.port_a_last_address = 29;
defparam ram_block5a0.port_a_logical_ram_depth = 30;
defparam ram_block5a0.port_a_logical_ram_width = 16;
defparam ram_block5a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a0.port_b_address_clear = "none";
defparam ram_block5a0.port_b_address_clock = "clock0";
defparam ram_block5a0.port_b_address_width = 5;
defparam ram_block5a0.port_b_data_out_clear = "clear0";
defparam ram_block5a0.port_b_data_out_clock = "clock0";
defparam ram_block5a0.port_b_data_width = 1;
defparam ram_block5a0.port_b_first_address = 0;
defparam ram_block5a0.port_b_first_bit_number = 0;
defparam ram_block5a0.port_b_last_address = 29;
defparam ram_block5a0.port_b_logical_ram_depth = 30;
defparam ram_block5a0.port_b_logical_ram_width = 16;
defparam ram_block5a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a0.port_b_read_enable_clock = "clock0";
defparam ram_block5a0.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a1_PORTBDATAOUT_bus));
defparam ram_block5a1.clk0_core_clock_enable = "ena0";
defparam ram_block5a1.clk0_input_clock_enable = "ena0";
defparam ram_block5a1.clk0_output_clock_enable = "ena0";
defparam ram_block5a1.data_interleave_offset_in_bits = 1;
defparam ram_block5a1.data_interleave_width_in_bits = 1;
defparam ram_block5a1.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|short_shift:short_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_euu:auto_generated|altsyncram_pbc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a1.mixed_port_feed_through_mode = "old";
defparam ram_block5a1.operation_mode = "dual_port";
defparam ram_block5a1.port_a_address_clear = "none";
defparam ram_block5a1.port_a_address_width = 5;
defparam ram_block5a1.port_a_data_out_clear = "none";
defparam ram_block5a1.port_a_data_out_clock = "none";
defparam ram_block5a1.port_a_data_width = 1;
defparam ram_block5a1.port_a_first_address = 0;
defparam ram_block5a1.port_a_first_bit_number = 1;
defparam ram_block5a1.port_a_last_address = 29;
defparam ram_block5a1.port_a_logical_ram_depth = 30;
defparam ram_block5a1.port_a_logical_ram_width = 16;
defparam ram_block5a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a1.port_b_address_clear = "none";
defparam ram_block5a1.port_b_address_clock = "clock0";
defparam ram_block5a1.port_b_address_width = 5;
defparam ram_block5a1.port_b_data_out_clear = "clear0";
defparam ram_block5a1.port_b_data_out_clock = "clock0";
defparam ram_block5a1.port_b_data_width = 1;
defparam ram_block5a1.port_b_first_address = 0;
defparam ram_block5a1.port_b_first_bit_number = 1;
defparam ram_block5a1.port_b_last_address = 29;
defparam ram_block5a1.port_b_logical_ram_depth = 30;
defparam ram_block5a1.port_b_logical_ram_width = 16;
defparam ram_block5a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a1.port_b_read_enable_clock = "clock0";
defparam ram_block5a1.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a2_PORTBDATAOUT_bus));
defparam ram_block5a2.clk0_core_clock_enable = "ena0";
defparam ram_block5a2.clk0_input_clock_enable = "ena0";
defparam ram_block5a2.clk0_output_clock_enable = "ena0";
defparam ram_block5a2.data_interleave_offset_in_bits = 1;
defparam ram_block5a2.data_interleave_width_in_bits = 1;
defparam ram_block5a2.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|short_shift:short_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_euu:auto_generated|altsyncram_pbc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a2.mixed_port_feed_through_mode = "old";
defparam ram_block5a2.operation_mode = "dual_port";
defparam ram_block5a2.port_a_address_clear = "none";
defparam ram_block5a2.port_a_address_width = 5;
defparam ram_block5a2.port_a_data_out_clear = "none";
defparam ram_block5a2.port_a_data_out_clock = "none";
defparam ram_block5a2.port_a_data_width = 1;
defparam ram_block5a2.port_a_first_address = 0;
defparam ram_block5a2.port_a_first_bit_number = 2;
defparam ram_block5a2.port_a_last_address = 29;
defparam ram_block5a2.port_a_logical_ram_depth = 30;
defparam ram_block5a2.port_a_logical_ram_width = 16;
defparam ram_block5a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a2.port_b_address_clear = "none";
defparam ram_block5a2.port_b_address_clock = "clock0";
defparam ram_block5a2.port_b_address_width = 5;
defparam ram_block5a2.port_b_data_out_clear = "clear0";
defparam ram_block5a2.port_b_data_out_clock = "clock0";
defparam ram_block5a2.port_b_data_width = 1;
defparam ram_block5a2.port_b_first_address = 0;
defparam ram_block5a2.port_b_first_bit_number = 2;
defparam ram_block5a2.port_b_last_address = 29;
defparam ram_block5a2.port_b_logical_ram_depth = 30;
defparam ram_block5a2.port_b_logical_ram_width = 16;
defparam ram_block5a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a2.port_b_read_enable_clock = "clock0";
defparam ram_block5a2.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a3_PORTBDATAOUT_bus));
defparam ram_block5a3.clk0_core_clock_enable = "ena0";
defparam ram_block5a3.clk0_input_clock_enable = "ena0";
defparam ram_block5a3.clk0_output_clock_enable = "ena0";
defparam ram_block5a3.data_interleave_offset_in_bits = 1;
defparam ram_block5a3.data_interleave_width_in_bits = 1;
defparam ram_block5a3.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|short_shift:short_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_euu:auto_generated|altsyncram_pbc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a3.mixed_port_feed_through_mode = "old";
defparam ram_block5a3.operation_mode = "dual_port";
defparam ram_block5a3.port_a_address_clear = "none";
defparam ram_block5a3.port_a_address_width = 5;
defparam ram_block5a3.port_a_data_out_clear = "none";
defparam ram_block5a3.port_a_data_out_clock = "none";
defparam ram_block5a3.port_a_data_width = 1;
defparam ram_block5a3.port_a_first_address = 0;
defparam ram_block5a3.port_a_first_bit_number = 3;
defparam ram_block5a3.port_a_last_address = 29;
defparam ram_block5a3.port_a_logical_ram_depth = 30;
defparam ram_block5a3.port_a_logical_ram_width = 16;
defparam ram_block5a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a3.port_b_address_clear = "none";
defparam ram_block5a3.port_b_address_clock = "clock0";
defparam ram_block5a3.port_b_address_width = 5;
defparam ram_block5a3.port_b_data_out_clear = "clear0";
defparam ram_block5a3.port_b_data_out_clock = "clock0";
defparam ram_block5a3.port_b_data_width = 1;
defparam ram_block5a3.port_b_first_address = 0;
defparam ram_block5a3.port_b_first_bit_number = 3;
defparam ram_block5a3.port_b_last_address = 29;
defparam ram_block5a3.port_b_logical_ram_depth = 30;
defparam ram_block5a3.port_b_logical_ram_width = 16;
defparam ram_block5a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a3.port_b_read_enable_clock = "clock0";
defparam ram_block5a3.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a4_PORTBDATAOUT_bus));
defparam ram_block5a4.clk0_core_clock_enable = "ena0";
defparam ram_block5a4.clk0_input_clock_enable = "ena0";
defparam ram_block5a4.clk0_output_clock_enable = "ena0";
defparam ram_block5a4.data_interleave_offset_in_bits = 1;
defparam ram_block5a4.data_interleave_width_in_bits = 1;
defparam ram_block5a4.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|short_shift:short_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_euu:auto_generated|altsyncram_pbc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a4.mixed_port_feed_through_mode = "old";
defparam ram_block5a4.operation_mode = "dual_port";
defparam ram_block5a4.port_a_address_clear = "none";
defparam ram_block5a4.port_a_address_width = 5;
defparam ram_block5a4.port_a_data_out_clear = "none";
defparam ram_block5a4.port_a_data_out_clock = "none";
defparam ram_block5a4.port_a_data_width = 1;
defparam ram_block5a4.port_a_first_address = 0;
defparam ram_block5a4.port_a_first_bit_number = 4;
defparam ram_block5a4.port_a_last_address = 29;
defparam ram_block5a4.port_a_logical_ram_depth = 30;
defparam ram_block5a4.port_a_logical_ram_width = 16;
defparam ram_block5a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a4.port_b_address_clear = "none";
defparam ram_block5a4.port_b_address_clock = "clock0";
defparam ram_block5a4.port_b_address_width = 5;
defparam ram_block5a4.port_b_data_out_clear = "clear0";
defparam ram_block5a4.port_b_data_out_clock = "clock0";
defparam ram_block5a4.port_b_data_width = 1;
defparam ram_block5a4.port_b_first_address = 0;
defparam ram_block5a4.port_b_first_bit_number = 4;
defparam ram_block5a4.port_b_last_address = 29;
defparam ram_block5a4.port_b_logical_ram_depth = 30;
defparam ram_block5a4.port_b_logical_ram_width = 16;
defparam ram_block5a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a4.port_b_read_enable_clock = "clock0";
defparam ram_block5a4.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a5_PORTBDATAOUT_bus));
defparam ram_block5a5.clk0_core_clock_enable = "ena0";
defparam ram_block5a5.clk0_input_clock_enable = "ena0";
defparam ram_block5a5.clk0_output_clock_enable = "ena0";
defparam ram_block5a5.data_interleave_offset_in_bits = 1;
defparam ram_block5a5.data_interleave_width_in_bits = 1;
defparam ram_block5a5.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|short_shift:short_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_euu:auto_generated|altsyncram_pbc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a5.mixed_port_feed_through_mode = "old";
defparam ram_block5a5.operation_mode = "dual_port";
defparam ram_block5a5.port_a_address_clear = "none";
defparam ram_block5a5.port_a_address_width = 5;
defparam ram_block5a5.port_a_data_out_clear = "none";
defparam ram_block5a5.port_a_data_out_clock = "none";
defparam ram_block5a5.port_a_data_width = 1;
defparam ram_block5a5.port_a_first_address = 0;
defparam ram_block5a5.port_a_first_bit_number = 5;
defparam ram_block5a5.port_a_last_address = 29;
defparam ram_block5a5.port_a_logical_ram_depth = 30;
defparam ram_block5a5.port_a_logical_ram_width = 16;
defparam ram_block5a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a5.port_b_address_clear = "none";
defparam ram_block5a5.port_b_address_clock = "clock0";
defparam ram_block5a5.port_b_address_width = 5;
defparam ram_block5a5.port_b_data_out_clear = "clear0";
defparam ram_block5a5.port_b_data_out_clock = "clock0";
defparam ram_block5a5.port_b_data_width = 1;
defparam ram_block5a5.port_b_first_address = 0;
defparam ram_block5a5.port_b_first_bit_number = 5;
defparam ram_block5a5.port_b_last_address = 29;
defparam ram_block5a5.port_b_logical_ram_depth = 30;
defparam ram_block5a5.port_b_logical_ram_width = 16;
defparam ram_block5a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a5.port_b_read_enable_clock = "clock0";
defparam ram_block5a5.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a6_PORTBDATAOUT_bus));
defparam ram_block5a6.clk0_core_clock_enable = "ena0";
defparam ram_block5a6.clk0_input_clock_enable = "ena0";
defparam ram_block5a6.clk0_output_clock_enable = "ena0";
defparam ram_block5a6.data_interleave_offset_in_bits = 1;
defparam ram_block5a6.data_interleave_width_in_bits = 1;
defparam ram_block5a6.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|short_shift:short_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_euu:auto_generated|altsyncram_pbc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a6.mixed_port_feed_through_mode = "old";
defparam ram_block5a6.operation_mode = "dual_port";
defparam ram_block5a6.port_a_address_clear = "none";
defparam ram_block5a6.port_a_address_width = 5;
defparam ram_block5a6.port_a_data_out_clear = "none";
defparam ram_block5a6.port_a_data_out_clock = "none";
defparam ram_block5a6.port_a_data_width = 1;
defparam ram_block5a6.port_a_first_address = 0;
defparam ram_block5a6.port_a_first_bit_number = 6;
defparam ram_block5a6.port_a_last_address = 29;
defparam ram_block5a6.port_a_logical_ram_depth = 30;
defparam ram_block5a6.port_a_logical_ram_width = 16;
defparam ram_block5a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a6.port_b_address_clear = "none";
defparam ram_block5a6.port_b_address_clock = "clock0";
defparam ram_block5a6.port_b_address_width = 5;
defparam ram_block5a6.port_b_data_out_clear = "clear0";
defparam ram_block5a6.port_b_data_out_clock = "clock0";
defparam ram_block5a6.port_b_data_width = 1;
defparam ram_block5a6.port_b_first_address = 0;
defparam ram_block5a6.port_b_first_bit_number = 6;
defparam ram_block5a6.port_b_last_address = 29;
defparam ram_block5a6.port_b_logical_ram_depth = 30;
defparam ram_block5a6.port_b_logical_ram_width = 16;
defparam ram_block5a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a6.port_b_read_enable_clock = "clock0";
defparam ram_block5a6.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a7_PORTBDATAOUT_bus));
defparam ram_block5a7.clk0_core_clock_enable = "ena0";
defparam ram_block5a7.clk0_input_clock_enable = "ena0";
defparam ram_block5a7.clk0_output_clock_enable = "ena0";
defparam ram_block5a7.data_interleave_offset_in_bits = 1;
defparam ram_block5a7.data_interleave_width_in_bits = 1;
defparam ram_block5a7.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|short_shift:short_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_euu:auto_generated|altsyncram_pbc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a7.mixed_port_feed_through_mode = "old";
defparam ram_block5a7.operation_mode = "dual_port";
defparam ram_block5a7.port_a_address_clear = "none";
defparam ram_block5a7.port_a_address_width = 5;
defparam ram_block5a7.port_a_data_out_clear = "none";
defparam ram_block5a7.port_a_data_out_clock = "none";
defparam ram_block5a7.port_a_data_width = 1;
defparam ram_block5a7.port_a_first_address = 0;
defparam ram_block5a7.port_a_first_bit_number = 7;
defparam ram_block5a7.port_a_last_address = 29;
defparam ram_block5a7.port_a_logical_ram_depth = 30;
defparam ram_block5a7.port_a_logical_ram_width = 16;
defparam ram_block5a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a7.port_b_address_clear = "none";
defparam ram_block5a7.port_b_address_clock = "clock0";
defparam ram_block5a7.port_b_address_width = 5;
defparam ram_block5a7.port_b_data_out_clear = "clear0";
defparam ram_block5a7.port_b_data_out_clock = "clock0";
defparam ram_block5a7.port_b_data_width = 1;
defparam ram_block5a7.port_b_first_address = 0;
defparam ram_block5a7.port_b_first_bit_number = 7;
defparam ram_block5a7.port_b_last_address = 29;
defparam ram_block5a7.port_b_logical_ram_depth = 30;
defparam ram_block5a7.port_b_logical_ram_width = 16;
defparam ram_block5a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a7.port_b_read_enable_clock = "clock0";
defparam ram_block5a7.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a8(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a8_PORTBDATAOUT_bus));
defparam ram_block5a8.clk0_core_clock_enable = "ena0";
defparam ram_block5a8.clk0_input_clock_enable = "ena0";
defparam ram_block5a8.clk0_output_clock_enable = "ena0";
defparam ram_block5a8.data_interleave_offset_in_bits = 1;
defparam ram_block5a8.data_interleave_width_in_bits = 1;
defparam ram_block5a8.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|short_shift:short_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_euu:auto_generated|altsyncram_pbc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a8.mixed_port_feed_through_mode = "old";
defparam ram_block5a8.operation_mode = "dual_port";
defparam ram_block5a8.port_a_address_clear = "none";
defparam ram_block5a8.port_a_address_width = 5;
defparam ram_block5a8.port_a_data_out_clear = "none";
defparam ram_block5a8.port_a_data_out_clock = "none";
defparam ram_block5a8.port_a_data_width = 1;
defparam ram_block5a8.port_a_first_address = 0;
defparam ram_block5a8.port_a_first_bit_number = 8;
defparam ram_block5a8.port_a_last_address = 29;
defparam ram_block5a8.port_a_logical_ram_depth = 30;
defparam ram_block5a8.port_a_logical_ram_width = 16;
defparam ram_block5a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a8.port_b_address_clear = "none";
defparam ram_block5a8.port_b_address_clock = "clock0";
defparam ram_block5a8.port_b_address_width = 5;
defparam ram_block5a8.port_b_data_out_clear = "clear0";
defparam ram_block5a8.port_b_data_out_clock = "clock0";
defparam ram_block5a8.port_b_data_width = 1;
defparam ram_block5a8.port_b_first_address = 0;
defparam ram_block5a8.port_b_first_bit_number = 8;
defparam ram_block5a8.port_b_last_address = 29;
defparam ram_block5a8.port_b_logical_ram_depth = 30;
defparam ram_block5a8.port_b_logical_ram_width = 16;
defparam ram_block5a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a8.port_b_read_enable_clock = "clock0";
defparam ram_block5a8.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a9(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a9_PORTBDATAOUT_bus));
defparam ram_block5a9.clk0_core_clock_enable = "ena0";
defparam ram_block5a9.clk0_input_clock_enable = "ena0";
defparam ram_block5a9.clk0_output_clock_enable = "ena0";
defparam ram_block5a9.data_interleave_offset_in_bits = 1;
defparam ram_block5a9.data_interleave_width_in_bits = 1;
defparam ram_block5a9.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|short_shift:short_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_euu:auto_generated|altsyncram_pbc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a9.mixed_port_feed_through_mode = "old";
defparam ram_block5a9.operation_mode = "dual_port";
defparam ram_block5a9.port_a_address_clear = "none";
defparam ram_block5a9.port_a_address_width = 5;
defparam ram_block5a9.port_a_data_out_clear = "none";
defparam ram_block5a9.port_a_data_out_clock = "none";
defparam ram_block5a9.port_a_data_width = 1;
defparam ram_block5a9.port_a_first_address = 0;
defparam ram_block5a9.port_a_first_bit_number = 9;
defparam ram_block5a9.port_a_last_address = 29;
defparam ram_block5a9.port_a_logical_ram_depth = 30;
defparam ram_block5a9.port_a_logical_ram_width = 16;
defparam ram_block5a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a9.port_b_address_clear = "none";
defparam ram_block5a9.port_b_address_clock = "clock0";
defparam ram_block5a9.port_b_address_width = 5;
defparam ram_block5a9.port_b_data_out_clear = "clear0";
defparam ram_block5a9.port_b_data_out_clock = "clock0";
defparam ram_block5a9.port_b_data_width = 1;
defparam ram_block5a9.port_b_first_address = 0;
defparam ram_block5a9.port_b_first_bit_number = 9;
defparam ram_block5a9.port_b_last_address = 29;
defparam ram_block5a9.port_b_logical_ram_depth = 30;
defparam ram_block5a9.port_b_logical_ram_width = 16;
defparam ram_block5a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a9.port_b_read_enable_clock = "clock0";
defparam ram_block5a9.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a10(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a10_PORTBDATAOUT_bus));
defparam ram_block5a10.clk0_core_clock_enable = "ena0";
defparam ram_block5a10.clk0_input_clock_enable = "ena0";
defparam ram_block5a10.clk0_output_clock_enable = "ena0";
defparam ram_block5a10.data_interleave_offset_in_bits = 1;
defparam ram_block5a10.data_interleave_width_in_bits = 1;
defparam ram_block5a10.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|short_shift:short_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_euu:auto_generated|altsyncram_pbc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a10.mixed_port_feed_through_mode = "old";
defparam ram_block5a10.operation_mode = "dual_port";
defparam ram_block5a10.port_a_address_clear = "none";
defparam ram_block5a10.port_a_address_width = 5;
defparam ram_block5a10.port_a_data_out_clear = "none";
defparam ram_block5a10.port_a_data_out_clock = "none";
defparam ram_block5a10.port_a_data_width = 1;
defparam ram_block5a10.port_a_first_address = 0;
defparam ram_block5a10.port_a_first_bit_number = 10;
defparam ram_block5a10.port_a_last_address = 29;
defparam ram_block5a10.port_a_logical_ram_depth = 30;
defparam ram_block5a10.port_a_logical_ram_width = 16;
defparam ram_block5a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a10.port_b_address_clear = "none";
defparam ram_block5a10.port_b_address_clock = "clock0";
defparam ram_block5a10.port_b_address_width = 5;
defparam ram_block5a10.port_b_data_out_clear = "clear0";
defparam ram_block5a10.port_b_data_out_clock = "clock0";
defparam ram_block5a10.port_b_data_width = 1;
defparam ram_block5a10.port_b_first_address = 0;
defparam ram_block5a10.port_b_first_bit_number = 10;
defparam ram_block5a10.port_b_last_address = 29;
defparam ram_block5a10.port_b_logical_ram_depth = 30;
defparam ram_block5a10.port_b_logical_ram_width = 16;
defparam ram_block5a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a10.port_b_read_enable_clock = "clock0";
defparam ram_block5a10.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a11(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a11_PORTBDATAOUT_bus));
defparam ram_block5a11.clk0_core_clock_enable = "ena0";
defparam ram_block5a11.clk0_input_clock_enable = "ena0";
defparam ram_block5a11.clk0_output_clock_enable = "ena0";
defparam ram_block5a11.data_interleave_offset_in_bits = 1;
defparam ram_block5a11.data_interleave_width_in_bits = 1;
defparam ram_block5a11.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|short_shift:short_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_euu:auto_generated|altsyncram_pbc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a11.mixed_port_feed_through_mode = "old";
defparam ram_block5a11.operation_mode = "dual_port";
defparam ram_block5a11.port_a_address_clear = "none";
defparam ram_block5a11.port_a_address_width = 5;
defparam ram_block5a11.port_a_data_out_clear = "none";
defparam ram_block5a11.port_a_data_out_clock = "none";
defparam ram_block5a11.port_a_data_width = 1;
defparam ram_block5a11.port_a_first_address = 0;
defparam ram_block5a11.port_a_first_bit_number = 11;
defparam ram_block5a11.port_a_last_address = 29;
defparam ram_block5a11.port_a_logical_ram_depth = 30;
defparam ram_block5a11.port_a_logical_ram_width = 16;
defparam ram_block5a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a11.port_b_address_clear = "none";
defparam ram_block5a11.port_b_address_clock = "clock0";
defparam ram_block5a11.port_b_address_width = 5;
defparam ram_block5a11.port_b_data_out_clear = "clear0";
defparam ram_block5a11.port_b_data_out_clock = "clock0";
defparam ram_block5a11.port_b_data_width = 1;
defparam ram_block5a11.port_b_first_address = 0;
defparam ram_block5a11.port_b_first_bit_number = 11;
defparam ram_block5a11.port_b_last_address = 29;
defparam ram_block5a11.port_b_logical_ram_depth = 30;
defparam ram_block5a11.port_b_logical_ram_width = 16;
defparam ram_block5a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a11.port_b_read_enable_clock = "clock0";
defparam ram_block5a11.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a12(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a12_PORTBDATAOUT_bus));
defparam ram_block5a12.clk0_core_clock_enable = "ena0";
defparam ram_block5a12.clk0_input_clock_enable = "ena0";
defparam ram_block5a12.clk0_output_clock_enable = "ena0";
defparam ram_block5a12.data_interleave_offset_in_bits = 1;
defparam ram_block5a12.data_interleave_width_in_bits = 1;
defparam ram_block5a12.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|short_shift:short_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_euu:auto_generated|altsyncram_pbc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a12.mixed_port_feed_through_mode = "old";
defparam ram_block5a12.operation_mode = "dual_port";
defparam ram_block5a12.port_a_address_clear = "none";
defparam ram_block5a12.port_a_address_width = 5;
defparam ram_block5a12.port_a_data_out_clear = "none";
defparam ram_block5a12.port_a_data_out_clock = "none";
defparam ram_block5a12.port_a_data_width = 1;
defparam ram_block5a12.port_a_first_address = 0;
defparam ram_block5a12.port_a_first_bit_number = 12;
defparam ram_block5a12.port_a_last_address = 29;
defparam ram_block5a12.port_a_logical_ram_depth = 30;
defparam ram_block5a12.port_a_logical_ram_width = 16;
defparam ram_block5a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a12.port_b_address_clear = "none";
defparam ram_block5a12.port_b_address_clock = "clock0";
defparam ram_block5a12.port_b_address_width = 5;
defparam ram_block5a12.port_b_data_out_clear = "clear0";
defparam ram_block5a12.port_b_data_out_clock = "clock0";
defparam ram_block5a12.port_b_data_width = 1;
defparam ram_block5a12.port_b_first_address = 0;
defparam ram_block5a12.port_b_first_bit_number = 12;
defparam ram_block5a12.port_b_last_address = 29;
defparam ram_block5a12.port_b_logical_ram_depth = 30;
defparam ram_block5a12.port_b_logical_ram_width = 16;
defparam ram_block5a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a12.port_b_read_enable_clock = "clock0";
defparam ram_block5a12.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a13(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a13_PORTBDATAOUT_bus));
defparam ram_block5a13.clk0_core_clock_enable = "ena0";
defparam ram_block5a13.clk0_input_clock_enable = "ena0";
defparam ram_block5a13.clk0_output_clock_enable = "ena0";
defparam ram_block5a13.data_interleave_offset_in_bits = 1;
defparam ram_block5a13.data_interleave_width_in_bits = 1;
defparam ram_block5a13.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|short_shift:short_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_euu:auto_generated|altsyncram_pbc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a13.mixed_port_feed_through_mode = "old";
defparam ram_block5a13.operation_mode = "dual_port";
defparam ram_block5a13.port_a_address_clear = "none";
defparam ram_block5a13.port_a_address_width = 5;
defparam ram_block5a13.port_a_data_out_clear = "none";
defparam ram_block5a13.port_a_data_out_clock = "none";
defparam ram_block5a13.port_a_data_width = 1;
defparam ram_block5a13.port_a_first_address = 0;
defparam ram_block5a13.port_a_first_bit_number = 13;
defparam ram_block5a13.port_a_last_address = 29;
defparam ram_block5a13.port_a_logical_ram_depth = 30;
defparam ram_block5a13.port_a_logical_ram_width = 16;
defparam ram_block5a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a13.port_b_address_clear = "none";
defparam ram_block5a13.port_b_address_clock = "clock0";
defparam ram_block5a13.port_b_address_width = 5;
defparam ram_block5a13.port_b_data_out_clear = "clear0";
defparam ram_block5a13.port_b_data_out_clock = "clock0";
defparam ram_block5a13.port_b_data_width = 1;
defparam ram_block5a13.port_b_first_address = 0;
defparam ram_block5a13.port_b_first_bit_number = 13;
defparam ram_block5a13.port_b_last_address = 29;
defparam ram_block5a13.port_b_logical_ram_depth = 30;
defparam ram_block5a13.port_b_logical_ram_width = 16;
defparam ram_block5a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a13.port_b_read_enable_clock = "clock0";
defparam ram_block5a13.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a14(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a14_PORTBDATAOUT_bus));
defparam ram_block5a14.clk0_core_clock_enable = "ena0";
defparam ram_block5a14.clk0_input_clock_enable = "ena0";
defparam ram_block5a14.clk0_output_clock_enable = "ena0";
defparam ram_block5a14.data_interleave_offset_in_bits = 1;
defparam ram_block5a14.data_interleave_width_in_bits = 1;
defparam ram_block5a14.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|short_shift:short_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_euu:auto_generated|altsyncram_pbc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a14.mixed_port_feed_through_mode = "old";
defparam ram_block5a14.operation_mode = "dual_port";
defparam ram_block5a14.port_a_address_clear = "none";
defparam ram_block5a14.port_a_address_width = 5;
defparam ram_block5a14.port_a_data_out_clear = "none";
defparam ram_block5a14.port_a_data_out_clock = "none";
defparam ram_block5a14.port_a_data_width = 1;
defparam ram_block5a14.port_a_first_address = 0;
defparam ram_block5a14.port_a_first_bit_number = 14;
defparam ram_block5a14.port_a_last_address = 29;
defparam ram_block5a14.port_a_logical_ram_depth = 30;
defparam ram_block5a14.port_a_logical_ram_width = 16;
defparam ram_block5a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a14.port_b_address_clear = "none";
defparam ram_block5a14.port_b_address_clock = "clock0";
defparam ram_block5a14.port_b_address_width = 5;
defparam ram_block5a14.port_b_data_out_clear = "clear0";
defparam ram_block5a14.port_b_data_out_clock = "clock0";
defparam ram_block5a14.port_b_data_width = 1;
defparam ram_block5a14.port_b_first_address = 0;
defparam ram_block5a14.port_b_first_bit_number = 14;
defparam ram_block5a14.port_b_last_address = 29;
defparam ram_block5a14.port_b_logical_ram_depth = 30;
defparam ram_block5a14.port_b_logical_ram_width = 16;
defparam ram_block5a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a14.port_b_read_enable_clock = "clock0";
defparam ram_block5a14.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block5a15(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block5a15_PORTBDATAOUT_bus));
defparam ram_block5a15.clk0_core_clock_enable = "ena0";
defparam ram_block5a15.clk0_input_clock_enable = "ena0";
defparam ram_block5a15.clk0_output_clock_enable = "ena0";
defparam ram_block5a15.data_interleave_offset_in_bits = 1;
defparam ram_block5a15.data_interleave_width_in_bits = 1;
defparam ram_block5a15.logical_ram_name = "packet_presence_detection:packet_presence_detection_0|dual_running_sum:running_sum_inst|short_shift:short_shift_inst|altshift_taps:ALTSHIFT_TAPS_component|shift_taps_euu:auto_generated|altsyncram_pbc1:altsyncram2|ALTSYNCRAM";
defparam ram_block5a15.mixed_port_feed_through_mode = "old";
defparam ram_block5a15.operation_mode = "dual_port";
defparam ram_block5a15.port_a_address_clear = "none";
defparam ram_block5a15.port_a_address_width = 5;
defparam ram_block5a15.port_a_data_out_clear = "none";
defparam ram_block5a15.port_a_data_out_clock = "none";
defparam ram_block5a15.port_a_data_width = 1;
defparam ram_block5a15.port_a_first_address = 0;
defparam ram_block5a15.port_a_first_bit_number = 15;
defparam ram_block5a15.port_a_last_address = 29;
defparam ram_block5a15.port_a_logical_ram_depth = 30;
defparam ram_block5a15.port_a_logical_ram_width = 16;
defparam ram_block5a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a15.port_b_address_clear = "none";
defparam ram_block5a15.port_b_address_clock = "clock0";
defparam ram_block5a15.port_b_address_width = 5;
defparam ram_block5a15.port_b_data_out_clear = "clear0";
defparam ram_block5a15.port_b_data_out_clock = "clock0";
defparam ram_block5a15.port_b_data_width = 1;
defparam ram_block5a15.port_b_first_address = 0;
defparam ram_block5a15.port_b_first_bit_number = 15;
defparam ram_block5a15.port_b_last_address = 29;
defparam ram_block5a15.port_b_logical_ram_depth = 30;
defparam ram_block5a15.port_b_logical_ram_width = 16;
defparam ram_block5a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block5a15.port_b_read_enable_clock = "clock0";
defparam ram_block5a15.ram_block_type = "M9K";

endmodule

module lms_dsp_cntr_5lg (
	counter_comb_bita41,
	always0,
	delay_reg_24_0,
	clock)/* synthesis synthesis_greybox=0 */;
output 	counter_comb_bita41;
input 	always0;
input 	delay_reg_24_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_reg_bit[4]~0_combout ;
wire \counter_reg_bit[0]~q ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_reg_bit[1]~q ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_reg_bit[2]~q ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_reg_bit[3]~q ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_reg_bit[4]~q ;
wire \counter_comb_bita4~COUT ;


fiftyfivenm_lcell_comb \counter_comb_bita4~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(counter_comb_bita41),
	.cout());
defparam \counter_comb_bita4~0 .lut_mask = 16'hF0F0;
defparam \counter_comb_bita4~0 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(\counter_reg_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5555;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter_reg_bit[4]~0 (
	.dataa(delay_reg_24_0),
	.datab(gnd),
	.datac(gnd),
	.datad(counter_comb_bita41),
	.cin(gnd),
	.combout(\counter_reg_bit[4]~0_combout ),
	.cout());
defparam \counter_reg_bit[4]~0 .lut_mask = 16'h00AA;
defparam \counter_reg_bit[4]~0 .sum_lutc_input = "datac";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!always0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\counter_reg_bit[4]~0_combout ),
	.q(\counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(\counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!always0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\counter_reg_bit[4]~0_combout ),
	.q(\counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(\counter_reg_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'hA50A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!always0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\counter_reg_bit[4]~0_combout ),
	.q(\counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(\counter_reg_bit[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!always0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\counter_reg_bit[4]~0_combout ),
	.q(\counter_reg_bit[3]~q ),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita4(
	.dataa(\counter_reg_bit[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'hA50A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!always0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\counter_reg_bit[4]~0_combout ),
	.q(\counter_reg_bit[4]~q ),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

endmodule

module lms_dsp_cntr_f5f (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	delay_reg_24_0,
	GND_port,
	clock)/* synthesis synthesis_greybox=0 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	delay_reg_24_0;
input 	GND_port;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \cmpr6|aneb_result_wire[0]~0_combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita4~0_combout ;
wire \cout_actual~combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita4~combout ;


lms_dsp_cmpr_hrb cmpr6(
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_4(counter_reg_bit_4),
	.aneb_result_wire_0(\cmpr6|aneb_result_wire[0]~0_combout ));

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\cout_actual~combout ),
	.ena(delay_reg_24_0),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\cout_actual~combout ),
	.ena(delay_reg_24_0),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\cout_actual~combout ),
	.ena(delay_reg_24_0),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\cout_actual~combout ),
	.ena(delay_reg_24_0),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\cout_actual~combout ),
	.ena(delay_reg_24_0),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'hA50A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'hA50A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter_comb_bita4~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita4~0_combout ),
	.cout());
defparam \counter_comb_bita4~0 .lut_mask = 16'hF0F0;
defparam \counter_comb_bita4~0 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb cout_actual(
	.dataa(\counter_comb_bita4~0_combout ),
	.datab(counter_reg_bit_0),
	.datac(\cmpr6|aneb_result_wire[0]~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\cout_actual~combout ),
	.cout());
defparam cout_actual.lut_mask = 16'hEAEA;
defparam cout_actual.sum_lutc_input = "datac";

endmodule

module lms_dsp_cmpr_hrb (
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	aneb_result_wire_0)/* synthesis synthesis_greybox=0 */;
input 	counter_reg_bit_1;
input 	counter_reg_bit_2;
input 	counter_reg_bit_3;
input 	counter_reg_bit_4;
output 	aneb_result_wire_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fiftyfivenm_lcell_comb \aneb_result_wire[0]~0 (
	.dataa(counter_reg_bit_2),
	.datab(counter_reg_bit_3),
	.datac(counter_reg_bit_4),
	.datad(counter_reg_bit_1),
	.cin(gnd),
	.combout(aneb_result_wire_0),
	.cout());
defparam \aneb_result_wire[0]~0 .lut_mask = 16'h0080;
defparam \aneb_result_wire[0]~0 .sum_lutc_input = "datac";

endmodule
